magic
tech gf180mcuD
magscale 1 10
timestamp 1751914308
<< nwell >>
rect -86 354 1430 870
<< pwell >>
rect -86 -86 1430 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 408 68 464 268
rect 568 68 624 268
rect 800 68 856 268
rect 960 68 1016 268
rect 1124 68 1180 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 528 440 584 716
rect 688 440 744 716
rect 800 440 856 716
rect 960 440 1016 716
rect 1124 440 1180 716
<< ndiff >>
rect 28 255 116 268
rect 28 209 41 255
rect 87 209 116 255
rect 28 68 116 209
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 68 408 268
rect 464 152 568 268
rect 464 106 493 152
rect 539 106 568 152
rect 464 68 568 106
rect 624 68 800 268
rect 856 127 960 268
rect 856 81 885 127
rect 931 81 960 127
rect 856 68 960 81
rect 1016 255 1124 268
rect 1016 209 1049 255
rect 1095 209 1124 255
rect 1016 68 1124 209
rect 1180 255 1300 268
rect 1180 81 1209 255
rect 1255 81 1300 255
rect 1180 68 1300 81
<< pdiff >>
rect 28 667 116 716
rect 28 453 41 667
rect 87 453 116 667
rect 28 440 116 453
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 440 528 716
rect 584 678 688 716
rect 584 632 613 678
rect 659 632 688 678
rect 584 440 688 632
rect 744 440 800 716
rect 856 703 960 716
rect 856 657 885 703
rect 931 657 960 703
rect 856 440 960 657
rect 1016 667 1124 716
rect 1016 453 1049 667
rect 1095 453 1124 667
rect 1016 440 1124 453
rect 1180 703 1300 716
rect 1180 453 1209 703
rect 1255 453 1300 703
rect 1180 440 1300 453
<< ndiffc >>
rect 41 209 87 255
rect 201 81 247 127
rect 493 106 539 152
rect 885 81 931 127
rect 1049 209 1095 255
rect 1209 81 1255 255
<< pdiffc >>
rect 41 453 87 667
rect 201 657 247 703
rect 613 632 659 678
rect 885 657 931 703
rect 1049 453 1095 667
rect 1209 453 1255 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 528 716 584 760
rect 688 716 744 760
rect 800 716 856 760
rect 960 716 1016 760
rect 1124 716 1180 760
rect 116 397 172 440
rect 276 397 332 440
rect 528 397 584 440
rect 688 397 744 440
rect 800 397 856 440
rect 960 397 1016 440
rect 116 376 200 397
rect 116 330 141 376
rect 187 330 200 376
rect 116 314 200 330
rect 276 377 360 397
rect 276 331 301 377
rect 347 331 360 377
rect 276 314 360 331
rect 408 376 480 397
rect 408 330 421 376
rect 467 330 480 376
rect 408 314 480 330
rect 528 380 601 397
rect 528 334 542 380
rect 588 351 601 380
rect 672 375 744 397
rect 588 334 624 351
rect 528 314 624 334
rect 672 329 685 375
rect 731 329 744 375
rect 672 314 744 329
rect 792 377 864 397
rect 792 331 805 377
rect 851 331 864 377
rect 792 314 864 331
rect 944 378 1016 397
rect 1124 378 1180 440
rect 944 332 957 378
rect 1003 332 1180 378
rect 944 314 1016 332
rect 116 268 172 314
rect 276 268 332 314
rect 408 268 464 314
rect 568 268 624 314
rect 800 268 856 314
rect 960 268 1016 314
rect 1124 268 1180 332
rect 116 24 172 68
rect 276 24 332 68
rect 408 24 464 68
rect 568 24 624 68
rect 800 24 856 68
rect 960 24 1016 68
rect 1124 24 1180 68
<< polycontact >>
rect 141 330 187 376
rect 301 331 347 377
rect 421 330 467 376
rect 542 334 588 380
rect 685 329 731 375
rect 805 331 851 377
rect 957 332 1003 378
<< metal1 >>
rect 0 724 1344 844
rect 201 703 247 724
rect 41 667 87 678
rect 885 703 931 724
rect 201 646 247 657
rect 544 632 613 678
rect 659 632 755 678
rect 1209 703 1255 724
rect 885 646 931 657
rect 1049 667 1115 678
rect 709 600 755 632
rect 87 554 497 600
rect 709 554 1003 600
rect 451 510 497 554
rect 41 255 87 453
rect 133 376 200 448
rect 133 330 141 376
rect 187 330 200 376
rect 133 314 200 330
rect 293 377 360 508
rect 451 464 588 510
rect 293 331 301 377
rect 347 331 360 377
rect 293 314 360 331
rect 421 376 467 388
rect 41 198 87 209
rect 141 245 187 314
rect 421 245 467 330
rect 542 380 588 464
rect 542 314 588 334
rect 672 375 744 508
rect 672 329 685 375
rect 731 329 744 375
rect 672 314 744 329
rect 792 377 864 508
rect 792 331 805 377
rect 851 331 864 377
rect 792 314 864 331
rect 957 378 1003 554
rect 685 245 731 314
rect 141 199 731 245
rect 957 230 1003 332
rect 793 184 1003 230
rect 1095 453 1115 667
rect 1049 255 1115 453
rect 1209 433 1255 453
rect 1095 209 1115 255
rect 1049 198 1115 209
rect 1209 255 1255 283
rect 793 152 839 184
rect 201 127 247 138
rect 441 106 493 152
rect 539 106 839 152
rect 885 127 931 138
rect 201 60 247 81
rect 885 60 931 81
rect 1209 60 1255 81
rect 0 -60 1344 60
<< labels >>
flabel metal1 s 0 724 1344 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1344 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 133 314 200 448 0 FreeSans 200 0 0 0 S
port 5 nsew signal input
flabel metal1 293 314 360 508 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 792 314 864 508 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
flabel metal1 672 314 744 508 0 FreeSans 200 0 0 0 S
port 5 nsew signal input
flabel metal1 1049 198 1115 678 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1344 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 1430 354
string MASKHINTS_PPLUS -86 354 1430 870
<< end >>
