magic
tech gf180mcuD
magscale 1 10
timestamp 1752061876
<< nwell >>
rect -86 354 1206 870
<< pwell >>
rect -86 -86 1206 354
<< nmos >>
rect 164 68 220 268
rect 452 68 508 268
rect 612 68 668 268
rect 772 68 828 268
rect 932 68 988 268
<< pmos >>
rect 164 440 220 716
rect 452 440 508 716
rect 612 440 668 716
rect 772 440 828 716
rect 932 440 988 716
<< ndiff >>
rect 75 244 164 268
rect 75 81 89 244
rect 135 81 164 244
rect 75 68 164 81
rect 220 255 308 268
rect 220 209 249 255
rect 295 209 308 255
rect 220 68 308 209
rect 364 127 452 268
rect 364 81 377 127
rect 423 81 452 127
rect 364 68 452 81
rect 508 244 612 268
rect 508 198 537 244
rect 583 198 612 244
rect 508 68 612 198
rect 668 127 772 268
rect 668 81 697 127
rect 743 81 772 127
rect 668 68 772 81
rect 828 255 932 268
rect 828 209 857 255
rect 903 209 932 255
rect 828 68 932 209
rect 988 127 1091 268
rect 988 81 1017 127
rect 1063 81 1091 127
rect 988 68 1091 81
<< pdiff >>
rect 75 703 164 716
rect 75 530 89 703
rect 135 530 164 703
rect 75 440 164 530
rect 220 667 308 716
rect 220 453 249 667
rect 295 453 308 667
rect 220 440 308 453
rect 364 597 452 716
rect 364 551 377 597
rect 423 551 452 597
rect 364 440 452 551
rect 508 703 612 716
rect 508 657 537 703
rect 583 657 612 703
rect 508 440 612 657
rect 668 678 772 716
rect 668 632 697 678
rect 743 632 772 678
rect 668 440 772 632
rect 828 569 932 716
rect 828 523 857 569
rect 903 523 932 569
rect 828 440 932 523
rect 988 678 1092 716
rect 988 632 1017 678
rect 1063 632 1092 678
rect 988 440 1092 632
<< ndiffc >>
rect 89 81 135 244
rect 249 209 295 255
rect 377 81 423 127
rect 537 198 583 244
rect 697 81 743 127
rect 857 209 903 255
rect 1017 81 1063 127
<< pdiffc >>
rect 89 530 135 703
rect 249 453 295 667
rect 377 551 423 597
rect 537 657 583 703
rect 697 632 743 678
rect 857 523 903 569
rect 1017 632 1063 678
<< polysilicon >>
rect 164 716 220 760
rect 452 716 508 760
rect 612 716 668 760
rect 772 716 828 760
rect 932 716 988 760
rect 164 395 220 440
rect 452 404 508 440
rect 612 404 668 440
rect 136 379 220 395
rect 136 333 149 379
rect 195 333 220 379
rect 136 320 220 333
rect 436 385 668 404
rect 772 403 828 440
rect 932 403 988 440
rect 436 339 449 385
rect 495 359 668 385
rect 495 339 508 359
rect 436 323 508 339
rect 164 268 220 320
rect 452 268 508 323
rect 612 268 668 359
rect 762 387 988 403
rect 762 341 775 387
rect 923 341 988 387
rect 762 322 988 341
rect 772 268 828 322
rect 932 268 988 322
rect 164 24 220 68
rect 452 24 508 68
rect 612 24 668 68
rect 772 24 828 68
rect 932 24 988 68
<< polycontact >>
rect 149 333 195 379
rect 449 339 495 385
rect 775 341 923 387
<< metal1 >>
rect 0 724 1120 844
rect 89 703 135 724
rect 537 703 583 724
rect 89 519 135 530
rect 249 667 295 678
rect 83 395 155 473
rect 537 646 583 657
rect 686 632 697 678
rect 743 632 1017 678
rect 1063 632 1074 678
rect 377 597 423 608
rect 686 585 732 632
rect 423 551 732 585
rect 969 569 1063 586
rect 377 539 732 551
rect 845 523 857 569
rect 903 523 1063 569
rect 83 379 195 395
rect 83 333 149 379
rect 83 309 195 333
rect 249 387 295 453
rect 436 387 500 404
rect 249 385 500 387
rect 249 341 449 385
rect 89 244 135 263
rect 249 255 295 341
rect 436 339 449 341
rect 495 339 500 385
rect 436 323 500 339
rect 666 387 923 403
rect 666 341 775 387
rect 666 322 923 341
rect 969 255 1063 523
rect 249 198 295 209
rect 537 244 857 255
rect 583 209 857 244
rect 903 209 1063 255
rect 537 187 583 198
rect 89 60 135 81
rect 377 127 423 138
rect 377 60 423 81
rect 697 127 743 138
rect 697 60 743 81
rect 1017 127 1063 138
rect 1017 60 1063 81
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 0 724 1120 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1120 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 969 210 1063 586 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 666 322 923 403 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 83 309 195 395 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
flabel metal1 83 395 155 473 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 1206 354
string MASKHINTS_PPLUS -86 354 1206 870
<< end >>
