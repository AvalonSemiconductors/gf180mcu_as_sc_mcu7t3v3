magic
tech gf180mcuD
magscale 1 10
timestamp 1753891287
<< nwell >>
rect -86 354 1654 870
<< pwell >>
rect -86 -86 1654 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 884 68 940 268
rect 1044 68 1100 268
rect 1204 68 1260 268
rect 1365 68 1421 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 884 440 940 716
rect 1044 440 1100 716
rect 1204 440 1260 716
rect 1365 440 1421 716
<< ndiff >>
rect 28 223 116 268
rect 28 177 41 223
rect 87 177 116 223
rect 28 68 116 177
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 213 436 268
rect 332 167 361 213
rect 407 167 436 213
rect 332 68 436 167
rect 492 244 596 268
rect 492 198 521 244
rect 567 198 596 244
rect 492 68 596 198
rect 652 152 740 268
rect 652 106 681 152
rect 727 106 740 152
rect 652 68 740 106
rect 796 152 884 268
rect 796 106 809 152
rect 855 106 884 152
rect 796 68 884 106
rect 940 244 1044 268
rect 940 198 969 244
rect 1015 198 1044 244
rect 940 68 1044 198
rect 1100 201 1204 268
rect 1100 155 1129 201
rect 1175 155 1204 201
rect 1100 68 1204 155
rect 1260 127 1365 268
rect 1260 81 1290 127
rect 1336 81 1365 127
rect 1260 68 1365 81
rect 1421 244 1509 268
rect 1421 198 1450 244
rect 1496 198 1509 244
rect 1421 68 1509 198
<< pdiff >>
rect 28 667 116 716
rect 28 453 41 667
rect 87 453 116 667
rect 28 440 116 453
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 667 436 716
rect 332 453 361 667
rect 407 453 436 667
rect 332 440 436 453
rect 492 703 596 716
rect 492 657 521 703
rect 567 657 596 703
rect 492 440 596 657
rect 652 667 884 716
rect 652 453 681 667
rect 727 453 782 667
rect 828 453 884 667
rect 652 440 884 453
rect 940 703 1044 716
rect 940 657 969 703
rect 1015 657 1044 703
rect 940 440 1044 657
rect 1100 667 1204 716
rect 1100 453 1129 667
rect 1175 453 1204 667
rect 1100 440 1204 453
rect 1260 510 1365 716
rect 1260 464 1290 510
rect 1336 464 1365 510
rect 1260 440 1365 464
rect 1421 667 1509 716
rect 1421 453 1450 667
rect 1496 453 1509 667
rect 1421 440 1509 453
<< ndiffc >>
rect 41 177 87 223
rect 201 81 247 127
rect 361 167 407 213
rect 521 198 567 244
rect 681 106 727 152
rect 809 106 855 152
rect 969 198 1015 244
rect 1129 155 1175 201
rect 1290 81 1336 127
rect 1450 198 1496 244
<< pdiffc >>
rect 41 453 87 667
rect 201 657 247 703
rect 361 453 407 667
rect 521 657 567 703
rect 681 453 727 667
rect 782 453 828 667
rect 969 657 1015 703
rect 1129 453 1175 667
rect 1290 464 1336 510
rect 1450 453 1496 667
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 884 716 940 760
rect 1044 716 1100 760
rect 1204 716 1260 760
rect 1365 716 1421 760
rect 116 391 172 440
rect 276 391 332 440
rect 116 378 332 391
rect 116 332 203 378
rect 249 332 332 378
rect 116 319 332 332
rect 116 268 172 319
rect 276 268 332 319
rect 436 391 492 440
rect 596 391 652 440
rect 436 378 652 391
rect 436 332 511 378
rect 557 332 652 378
rect 436 319 652 332
rect 436 268 492 319
rect 596 268 652 319
rect 884 391 940 440
rect 1044 391 1100 440
rect 1204 391 1260 440
rect 1365 391 1421 440
rect 884 378 1100 391
rect 884 332 1011 378
rect 1057 332 1100 378
rect 884 319 1100 332
rect 1182 378 1421 391
rect 1182 332 1219 378
rect 1265 332 1421 378
rect 1182 319 1421 332
rect 884 268 940 319
rect 1044 268 1100 319
rect 1204 268 1260 319
rect 1365 268 1421 319
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 884 24 940 68
rect 1044 24 1100 68
rect 1204 24 1260 68
rect 1365 24 1421 68
<< polycontact >>
rect 203 332 249 378
rect 511 332 557 378
rect 1011 332 1057 378
rect 1219 332 1265 378
<< metal1 >>
rect 0 724 1568 844
rect 201 703 247 724
rect 41 667 87 678
rect 521 703 567 724
rect 201 646 247 657
rect 361 667 407 678
rect 87 544 361 590
rect 41 440 87 453
rect 969 703 1015 724
rect 521 646 567 657
rect 681 667 727 678
rect 407 544 681 590
rect 361 440 407 453
rect 782 667 828 678
rect 727 544 782 590
rect 681 440 727 453
rect 969 646 1015 657
rect 1129 667 1496 678
rect 828 544 1129 590
rect 782 440 828 453
rect 1175 632 1450 667
rect 1271 464 1290 510
rect 1336 464 1403 510
rect 1129 440 1175 453
rect 116 378 332 385
rect 116 332 203 378
rect 249 332 332 378
rect 116 326 332 332
rect 436 378 652 385
rect 436 332 511 378
rect 557 332 652 378
rect 436 326 652 332
rect 884 378 1100 385
rect 884 332 1011 378
rect 1057 332 1100 378
rect 884 326 1100 332
rect 1182 378 1300 385
rect 1182 332 1219 378
rect 1265 332 1300 378
rect 1182 326 1300 332
rect 1346 244 1403 464
rect 1450 440 1496 453
rect 41 230 87 234
rect 41 223 407 230
rect 87 213 407 223
rect 87 184 361 213
rect 41 160 87 177
rect 494 198 521 244
rect 567 198 969 244
rect 1015 198 1026 244
rect 1129 201 1450 244
rect 361 152 407 167
rect 1175 198 1450 201
rect 1496 198 1507 244
rect 1129 152 1175 155
rect 201 127 247 138
rect 361 106 681 152
rect 727 106 739 152
rect 794 106 809 152
rect 855 106 1175 152
rect 1290 127 1336 138
rect 201 60 247 81
rect 1290 60 1336 81
rect 0 -60 1568 60
<< labels >>
flabel metal1 s 0 724 1568 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1568 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 116 326 332 385 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 436 326 652 385 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 884 326 1100 385 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 1346 198 1403 510 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel metal1 1182 326 1300 385 0 FreeSans 200 0 0 0 D
port 9 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 1654 354
string MASKHINTS_PPLUS -86 354 1654 870
<< end >>
