magic
tech gf180mcuD
magscale 1 10
timestamp 1751559330
<< nwell >>
rect -86 354 2102 870
<< pwell >>
rect -86 -86 2102 354
<< nmos >>
rect 116 68 172 212
rect 276 68 332 212
rect 436 68 492 212
rect 596 68 652 212
rect 756 68 812 212
rect 916 68 972 212
rect 1076 68 1132 212
rect 1236 68 1292 212
rect 1396 68 1452 212
rect 1556 68 1612 212
rect 1716 68 1772 212
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1396 440 1452 716
rect 1556 440 1612 716
rect 1716 440 1772 716
<< ndiff >>
rect 28 132 116 212
rect 28 86 41 132
rect 87 86 116 132
rect 28 68 116 86
rect 172 199 276 212
rect 172 153 201 199
rect 247 153 276 199
rect 172 68 276 153
rect 332 129 436 212
rect 332 83 361 129
rect 407 83 436 129
rect 332 68 436 83
rect 492 199 596 212
rect 492 153 521 199
rect 567 153 596 199
rect 492 68 596 153
rect 652 127 756 212
rect 652 81 681 127
rect 727 81 756 127
rect 652 68 756 81
rect 812 199 916 212
rect 812 153 841 199
rect 887 153 916 199
rect 812 68 916 153
rect 972 127 1076 212
rect 972 81 1001 127
rect 1047 81 1076 127
rect 972 68 1076 81
rect 1132 199 1236 212
rect 1132 153 1161 199
rect 1207 153 1236 199
rect 1132 68 1236 153
rect 1292 127 1396 212
rect 1292 81 1321 127
rect 1367 81 1396 127
rect 1292 68 1396 81
rect 1452 199 1556 212
rect 1452 153 1481 199
rect 1527 153 1556 199
rect 1452 68 1556 153
rect 1612 127 1716 212
rect 1612 81 1641 127
rect 1687 81 1716 127
rect 1612 68 1716 81
rect 1772 199 1988 212
rect 1772 153 1801 199
rect 1847 153 1988 199
rect 1772 68 1988 153
<< pdiff >>
rect 28 694 116 716
rect 28 648 41 694
rect 87 648 116 694
rect 28 440 116 648
rect 172 667 276 716
rect 172 453 201 667
rect 247 453 276 667
rect 172 440 276 453
rect 332 694 436 716
rect 332 464 361 694
rect 407 464 436 694
rect 332 440 436 464
rect 492 667 596 716
rect 492 453 521 667
rect 567 453 596 667
rect 492 440 596 453
rect 652 696 756 716
rect 652 453 681 696
rect 727 453 756 696
rect 652 440 756 453
rect 812 667 916 716
rect 812 453 841 667
rect 887 453 916 667
rect 812 440 916 453
rect 972 703 1076 716
rect 972 453 1001 703
rect 1047 453 1076 703
rect 972 440 1076 453
rect 1132 667 1236 716
rect 1132 453 1161 667
rect 1207 453 1236 667
rect 1132 440 1236 453
rect 1292 703 1396 716
rect 1292 453 1321 703
rect 1367 453 1396 703
rect 1292 440 1396 453
rect 1452 667 1556 716
rect 1452 453 1481 667
rect 1527 453 1556 667
rect 1452 440 1556 453
rect 1612 703 1716 716
rect 1612 453 1641 703
rect 1687 453 1716 703
rect 1612 440 1716 453
rect 1772 667 1988 716
rect 1772 453 1801 667
rect 1847 453 1988 667
rect 1772 440 1988 453
<< ndiffc >>
rect 41 86 87 132
rect 201 153 247 199
rect 361 83 407 129
rect 521 153 567 199
rect 681 81 727 127
rect 841 153 887 199
rect 1001 81 1047 127
rect 1161 153 1207 199
rect 1321 81 1367 127
rect 1481 153 1527 199
rect 1641 81 1687 127
rect 1801 153 1847 199
<< pdiffc >>
rect 41 648 87 694
rect 201 453 247 667
rect 361 464 407 694
rect 521 453 567 667
rect 681 453 727 696
rect 841 453 887 667
rect 1001 453 1047 703
rect 1161 453 1207 667
rect 1321 453 1367 703
rect 1481 453 1527 667
rect 1641 453 1687 703
rect 1801 453 1847 667
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1396 716 1452 760
rect 1556 716 1612 761
rect 1716 716 1772 761
rect 116 412 172 440
rect 276 412 332 440
rect 74 393 332 412
rect 436 393 492 440
rect 596 399 652 440
rect 756 399 812 440
rect 74 389 492 393
rect 74 343 95 389
rect 141 345 492 389
rect 141 343 332 345
rect 74 322 332 343
rect 116 212 172 322
rect 276 212 332 322
rect 436 212 492 345
rect 544 382 812 399
rect 544 336 557 382
rect 784 378 812 382
rect 916 378 972 440
rect 1076 378 1132 440
rect 1236 378 1292 440
rect 1396 378 1452 440
rect 1556 378 1612 440
rect 1716 378 1772 440
rect 784 336 1772 378
rect 544 332 1772 336
rect 544 322 812 332
rect 596 212 652 322
rect 756 212 812 322
rect 916 212 972 332
rect 1076 212 1132 332
rect 1236 212 1292 332
rect 1396 212 1452 332
rect 1556 212 1612 332
rect 1716 212 1772 332
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1396 24 1452 68
rect 1556 24 1612 68
rect 1716 24 1772 68
<< polycontact >>
rect 95 343 141 389
rect 557 336 784 382
<< metal1 >>
rect 0 724 2016 844
rect 41 694 87 724
rect 361 694 407 724
rect 41 637 87 648
rect 201 667 247 678
rect 41 412 117 481
rect 681 696 727 724
rect 361 453 407 464
rect 521 667 567 678
rect 41 389 154 412
rect 41 343 95 389
rect 141 343 154 389
rect 41 322 154 343
rect 201 407 247 453
rect 521 407 567 453
rect 1001 703 1047 724
rect 681 436 727 453
rect 841 667 887 678
rect 201 399 567 407
rect 201 387 613 399
rect 841 396 887 453
rect 1321 703 1367 724
rect 1001 442 1047 453
rect 1161 667 1207 678
rect 1161 396 1207 453
rect 1641 703 1687 724
rect 1321 442 1367 453
rect 1481 667 1527 678
rect 1481 396 1527 453
rect 1641 442 1687 453
rect 1801 667 1847 678
rect 1801 396 1847 453
rect 201 382 795 387
rect 201 361 557 382
rect 41 291 117 322
rect 201 199 247 361
rect 41 132 87 147
rect 201 142 247 153
rect 521 336 557 361
rect 784 336 795 382
rect 521 332 795 336
rect 521 322 613 332
rect 521 199 567 322
rect 841 314 1847 396
rect 841 199 887 314
rect 521 142 567 153
rect 41 60 87 86
rect 361 129 407 140
rect 361 60 407 83
rect 681 127 727 159
rect 1161 199 1207 314
rect 1481 199 1527 314
rect 841 142 887 153
rect 681 60 727 81
rect 1001 127 1047 153
rect 1161 142 1207 153
rect 1001 60 1047 81
rect 1321 127 1367 153
rect 1481 142 1527 153
rect 1801 199 1847 314
rect 1321 60 1367 81
rect 1641 127 1687 150
rect 1801 142 1847 153
rect 1641 60 1687 81
rect 0 -60 2016 60
<< labels >>
flabel metal1 s 0 724 2016 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2016 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 41 322 154 412 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 841 314 1847 396 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2016 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
