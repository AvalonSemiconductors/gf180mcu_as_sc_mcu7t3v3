magic
tech gf180mcuD
magscale 1 10
timestamp 1759840351
<< nwell >>
rect -86 354 2326 870
<< pwell >>
rect -86 -86 2326 354
<< nmos >>
rect 164 68 220 268
rect 452 68 508 268
rect 612 68 668 268
rect 772 68 828 268
rect 932 68 988 268
rect 1092 68 1148 268
rect 1252 68 1308 268
rect 1540 68 1596 268
rect 1700 68 1756 268
rect 1860 68 1916 268
rect 2020 68 2076 268
<< pmos >>
rect 164 440 220 716
rect 452 440 508 716
rect 612 440 668 716
rect 772 440 828 716
rect 932 440 988 716
rect 1092 440 1148 716
rect 1252 440 1308 716
rect 1540 440 1596 716
rect 1700 440 1756 716
rect 1860 440 1916 716
rect 2020 440 2076 716
<< ndiff >>
rect 70 127 164 268
rect 70 81 83 127
rect 129 81 164 127
rect 70 68 164 81
rect 220 255 308 268
rect 220 209 249 255
rect 295 209 308 255
rect 220 68 308 209
rect 364 127 452 268
rect 364 81 377 127
rect 423 81 452 127
rect 364 68 452 81
rect 508 68 612 268
rect 668 251 772 268
rect 668 205 697 251
rect 743 205 772 251
rect 668 68 772 205
rect 828 68 932 268
rect 988 127 1092 268
rect 988 81 1017 127
rect 1063 81 1092 127
rect 988 68 1092 81
rect 1148 251 1252 268
rect 1148 205 1177 251
rect 1223 205 1252 251
rect 1148 68 1252 205
rect 1308 127 1540 268
rect 1308 81 1337 127
rect 1510 81 1540 127
rect 1308 68 1540 81
rect 1596 255 1700 268
rect 1596 209 1625 255
rect 1671 209 1700 255
rect 1596 68 1700 209
rect 1756 127 1860 268
rect 1756 81 1785 127
rect 1831 81 1860 127
rect 1756 68 1860 81
rect 1916 255 2020 268
rect 1916 209 1945 255
rect 1991 209 2020 255
rect 1916 68 2020 209
rect 2076 127 2182 268
rect 2076 81 2105 127
rect 2151 81 2182 127
rect 2076 68 2182 81
<< pdiff >>
rect 72 703 164 716
rect 72 514 85 703
rect 131 514 164 703
rect 72 440 164 514
rect 220 667 308 716
rect 220 453 249 667
rect 295 453 308 667
rect 220 440 308 453
rect 364 600 452 716
rect 364 554 377 600
rect 423 554 452 600
rect 364 440 452 554
rect 508 703 612 716
rect 508 657 537 703
rect 583 657 612 703
rect 508 440 612 657
rect 668 600 772 716
rect 668 554 697 600
rect 743 554 772 600
rect 668 440 772 554
rect 828 703 932 716
rect 828 657 857 703
rect 903 657 932 703
rect 828 440 932 657
rect 988 639 1092 716
rect 988 593 1017 639
rect 1063 593 1092 639
rect 988 440 1092 593
rect 1148 499 1252 716
rect 1148 453 1177 499
rect 1223 453 1252 499
rect 1148 440 1252 453
rect 1308 652 1396 716
rect 1308 606 1337 652
rect 1383 606 1396 652
rect 1308 440 1396 606
rect 1452 703 1540 716
rect 1452 657 1465 703
rect 1511 657 1540 703
rect 1452 440 1540 657
rect 1596 667 1700 716
rect 1596 453 1625 667
rect 1671 453 1700 667
rect 1596 440 1700 453
rect 1756 703 1860 716
rect 1756 657 1785 703
rect 1831 657 1860 703
rect 1756 440 1860 657
rect 1916 667 2020 716
rect 1916 453 1945 667
rect 1991 453 2020 667
rect 1916 440 2020 453
rect 2076 703 2182 716
rect 2076 657 2105 703
rect 2151 657 2182 703
rect 2076 440 2182 657
<< ndiffc >>
rect 83 81 129 127
rect 249 209 295 255
rect 377 81 423 127
rect 697 205 743 251
rect 1017 81 1063 127
rect 1177 205 1223 251
rect 1337 81 1510 127
rect 1625 209 1671 255
rect 1785 81 1831 127
rect 1945 209 1991 255
rect 2105 81 2151 127
<< pdiffc >>
rect 85 514 131 703
rect 249 453 295 667
rect 377 554 423 600
rect 537 657 583 703
rect 697 554 743 600
rect 857 657 903 703
rect 1017 593 1063 639
rect 1177 453 1223 499
rect 1337 606 1383 652
rect 1465 657 1511 703
rect 1625 453 1671 667
rect 1785 657 1831 703
rect 1945 453 1991 667
rect 2105 657 2151 703
<< polysilicon >>
rect 164 716 220 760
rect 452 716 508 760
rect 612 716 668 760
rect 772 716 828 760
rect 932 716 988 760
rect 1092 716 1148 760
rect 1252 716 1308 760
rect 1540 716 1596 760
rect 1700 716 1756 760
rect 1860 716 1916 760
rect 2020 716 2076 760
rect 164 391 220 440
rect 131 378 220 391
rect 452 390 508 440
rect 131 332 144 378
rect 190 332 220 378
rect 131 319 220 332
rect 164 268 220 319
rect 427 377 508 390
rect 427 331 443 377
rect 489 331 508 377
rect 427 318 508 331
rect 452 268 508 318
rect 612 390 668 440
rect 772 390 828 440
rect 612 377 828 390
rect 932 386 988 440
rect 612 331 625 377
rect 815 331 828 377
rect 612 318 828 331
rect 612 268 668 318
rect 772 268 828 318
rect 908 373 989 386
rect 908 327 926 373
rect 972 327 989 373
rect 908 314 989 327
rect 1092 373 1148 440
rect 1252 392 1308 440
rect 1252 375 1361 392
rect 1540 389 1596 440
rect 1252 373 1300 375
rect 1092 329 1300 373
rect 1346 329 1361 375
rect 1092 327 1361 329
rect 932 268 988 314
rect 1092 268 1148 327
rect 1252 313 1361 327
rect 1497 377 1596 389
rect 1700 377 1756 440
rect 1860 377 1916 440
rect 2020 377 2076 440
rect 1497 372 2076 377
rect 1497 326 1514 372
rect 1560 326 2076 372
rect 1497 324 2076 326
rect 1252 268 1308 313
rect 1497 309 1596 324
rect 1540 268 1596 309
rect 1700 268 1756 324
rect 1860 268 1916 324
rect 2020 268 2076 324
rect 164 24 220 68
rect 452 24 508 68
rect 612 24 668 68
rect 772 24 828 68
rect 932 24 988 68
rect 1092 24 1148 68
rect 1252 24 1308 68
rect 1540 24 1596 68
rect 1700 24 1756 68
rect 1860 24 1916 68
rect 2020 24 2076 68
<< polycontact >>
rect 144 332 190 378
rect 443 331 489 377
rect 625 331 815 377
rect 926 327 972 373
rect 1300 329 1346 375
rect 1514 326 1560 372
<< metal1 >>
rect 0 724 2240 844
rect 85 703 131 724
rect 537 703 583 724
rect 85 503 131 514
rect 249 667 295 678
rect 122 378 203 457
rect 122 332 144 378
rect 190 332 203 378
rect 122 296 203 332
rect 537 646 583 657
rect 857 703 903 724
rect 1465 703 1511 724
rect 857 646 903 657
rect 1017 652 1383 678
rect 1017 639 1337 652
rect 377 600 423 616
rect 423 554 697 600
rect 743 593 1017 600
rect 1063 632 1337 639
rect 1785 703 1831 724
rect 1465 646 1511 657
rect 1622 667 1675 678
rect 1337 594 1383 606
rect 743 554 1063 593
rect 377 539 423 554
rect 249 389 295 453
rect 465 462 954 508
rect 465 391 511 462
rect 427 389 511 391
rect 249 377 511 389
rect 249 331 443 377
rect 489 331 511 377
rect 249 319 511 331
rect 249 255 295 319
rect 427 318 511 319
rect 612 377 828 390
rect 612 331 625 377
rect 815 331 828 377
rect 612 318 828 331
rect 908 386 954 462
rect 1165 499 1223 524
rect 1165 453 1177 499
rect 908 373 989 386
rect 908 327 926 373
rect 972 327 989 373
rect 908 314 989 327
rect 1165 251 1223 453
rect 1283 375 1361 462
rect 1622 453 1625 667
rect 1671 453 1675 667
rect 2105 703 2151 724
rect 1785 646 1831 657
rect 1940 667 1993 678
rect 1283 329 1300 375
rect 1346 329 1361 375
rect 1283 313 1361 329
rect 1497 372 1574 389
rect 1497 326 1514 372
rect 1560 326 1574 372
rect 1497 309 1574 326
rect 1622 379 1675 453
rect 1940 453 1945 667
rect 1991 453 1993 667
rect 2105 646 2151 657
rect 1940 379 1993 453
rect 1622 329 1993 379
rect 1497 251 1543 309
rect 249 197 295 209
rect 672 205 697 251
rect 743 205 1177 251
rect 1223 205 1543 251
rect 1622 255 1675 329
rect 1622 209 1625 255
rect 1671 209 1675 255
rect 1622 198 1675 209
rect 1940 255 1993 329
rect 1940 209 1945 255
rect 1991 209 1993 255
rect 1940 198 1993 209
rect 83 127 129 138
rect 83 60 129 81
rect 377 127 423 138
rect 377 60 423 81
rect 1017 127 1063 138
rect 1017 60 1063 81
rect 1337 127 1510 138
rect 1337 60 1510 81
rect 1785 127 1831 138
rect 1785 60 1831 81
rect 2105 127 2151 138
rect 2105 60 2151 81
rect 0 -60 2240 60
<< labels >>
flabel metal1 s 0 724 2240 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2240 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 1283 313 1361 462 0 FreeSans 200 0 0 0 C
port 6 nsew signal input
flabel metal1 612 318 828 390 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 122 296 203 457 0 FreeSans 200 0 0 0 A
port 8 nsew signal input
flabel metal1 1622 198 1675 678 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 1940 198 1993 678 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2240 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 2256 354
string MASKHINTS_PPLUS -16 354 2256 830
<< end >>
