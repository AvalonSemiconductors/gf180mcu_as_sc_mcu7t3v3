magic
tech gf180mcuD
magscale 1 10
timestamp 1753869255
<< nwell >>
rect -86 354 1654 870
<< pwell >>
rect -86 -86 1654 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 564 68 620 268
rect 724 68 780 268
rect 884 68 940 268
rect 1044 68 1100 268
rect 1204 68 1260 268
rect 1364 68 1420 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 564 440 620 716
rect 724 440 780 716
rect 884 440 940 716
rect 1044 440 1100 716
rect 1204 440 1260 716
rect 1364 440 1420 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 68 276 268
rect 332 152 420 268
rect 332 106 361 152
rect 407 106 420 152
rect 332 68 420 106
rect 476 152 564 268
rect 476 106 489 152
rect 535 106 564 152
rect 476 68 564 106
rect 620 68 724 268
rect 780 127 884 268
rect 780 81 809 127
rect 855 81 884 127
rect 780 68 884 81
rect 940 255 1044 268
rect 940 209 969 255
rect 1015 209 1044 255
rect 940 68 1044 209
rect 1100 255 1204 268
rect 1100 81 1129 255
rect 1175 81 1204 255
rect 1100 68 1204 81
rect 1260 254 1364 268
rect 1260 208 1289 254
rect 1335 208 1364 254
rect 1260 68 1364 208
rect 1420 255 1508 268
rect 1420 81 1449 255
rect 1495 81 1508 255
rect 1420 68 1508 81
<< pdiff >>
rect 28 667 116 716
rect 28 459 41 667
rect 87 459 116 667
rect 28 440 116 459
rect 172 586 276 716
rect 172 540 201 586
rect 247 540 276 586
rect 172 440 276 540
rect 332 678 420 716
rect 332 632 361 678
rect 407 632 420 678
rect 332 440 420 632
rect 476 703 564 716
rect 476 657 489 703
rect 535 657 564 703
rect 476 440 564 657
rect 620 611 724 716
rect 620 565 649 611
rect 695 565 724 611
rect 620 440 724 565
rect 780 703 884 716
rect 780 657 809 703
rect 855 657 884 703
rect 780 440 884 657
rect 940 667 1044 716
rect 940 453 969 667
rect 1015 453 1044 667
rect 940 440 1044 453
rect 1100 703 1204 716
rect 1100 453 1129 703
rect 1175 453 1204 703
rect 1100 440 1204 453
rect 1260 667 1364 716
rect 1260 453 1289 667
rect 1335 453 1364 667
rect 1260 440 1364 453
rect 1420 703 1508 716
rect 1420 453 1449 703
rect 1495 453 1508 703
rect 1420 440 1508 453
<< ndiffc >>
rect 41 81 87 127
rect 361 106 407 152
rect 489 106 535 152
rect 809 81 855 127
rect 969 209 1015 255
rect 1129 81 1175 255
rect 1289 208 1335 254
rect 1449 81 1495 255
<< pdiffc >>
rect 41 459 87 667
rect 201 540 247 586
rect 361 632 407 678
rect 489 657 535 703
rect 649 565 695 611
rect 809 657 855 703
rect 969 453 1015 667
rect 1129 453 1175 703
rect 1289 453 1335 667
rect 1449 453 1495 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 564 716 620 760
rect 724 716 780 760
rect 884 716 940 760
rect 1044 716 1100 760
rect 1204 716 1260 760
rect 1364 716 1420 760
rect 116 394 172 440
rect 276 402 332 440
rect 564 402 620 440
rect 724 402 780 440
rect 70 379 172 394
rect 70 333 98 379
rect 144 333 172 379
rect 70 318 172 333
rect 116 268 172 318
rect 253 376 358 402
rect 253 330 282 376
rect 328 330 358 376
rect 253 312 358 330
rect 478 371 620 402
rect 478 325 492 371
rect 538 325 620 371
rect 478 312 620 325
rect 699 378 804 402
rect 884 389 940 440
rect 699 332 729 378
rect 775 332 804 378
rect 699 312 804 332
rect 859 376 940 389
rect 1044 376 1100 440
rect 1204 376 1260 440
rect 1364 376 1420 440
rect 859 330 872 376
rect 918 330 1420 376
rect 859 317 940 330
rect 276 268 332 312
rect 564 268 620 312
rect 724 268 780 312
rect 884 268 940 317
rect 1044 268 1100 330
rect 1204 268 1260 330
rect 1364 268 1420 330
rect 116 24 172 68
rect 276 24 332 68
rect 564 24 620 68
rect 724 24 780 68
rect 884 24 940 68
rect 1044 24 1100 68
rect 1204 24 1260 68
rect 1364 24 1420 68
<< polycontact >>
rect 98 333 144 379
rect 282 330 328 376
rect 492 325 538 371
rect 729 332 775 378
rect 872 330 918 376
<< metal1 >>
rect 0 724 1568 844
rect 489 703 535 724
rect 41 667 361 678
rect 87 632 361 667
rect 407 632 418 678
rect 489 646 535 657
rect 809 703 855 724
rect 1129 703 1175 724
rect 809 646 855 657
rect 969 667 1036 678
rect 649 611 695 632
rect 180 540 201 586
rect 247 565 649 586
rect 247 540 695 565
rect 87 459 918 494
rect 41 448 918 459
rect 67 379 172 402
rect 67 333 98 379
rect 144 333 172 379
rect 67 312 172 333
rect 253 376 358 402
rect 253 330 282 376
rect 328 330 358 376
rect 253 312 358 330
rect 478 371 583 402
rect 478 325 492 371
rect 538 325 583 371
rect 478 312 583 325
rect 699 378 804 402
rect 699 332 729 378
rect 775 332 804 378
rect 699 312 804 332
rect 872 376 918 448
rect 872 249 918 330
rect 650 203 918 249
rect 1015 453 1036 667
rect 969 376 1036 453
rect 1449 703 1495 724
rect 1129 431 1175 453
rect 1289 667 1356 678
rect 1335 453 1356 667
rect 1289 376 1356 453
rect 1449 431 1495 453
rect 969 330 1356 376
rect 969 255 1036 330
rect 1015 209 1036 255
rect 650 152 696 203
rect 969 196 1036 209
rect 1129 255 1175 277
rect 41 127 87 138
rect 327 106 361 152
rect 407 106 489 152
rect 535 106 696 152
rect 809 127 855 138
rect 41 60 87 81
rect 809 60 855 81
rect 1289 254 1356 330
rect 1335 208 1356 254
rect 1289 196 1356 208
rect 1449 255 1495 277
rect 1129 60 1175 81
rect 1449 60 1495 81
rect 0 -60 1568 60
<< labels >>
flabel metal1 s 0 724 1568 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1568 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 67 312 172 402 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 253 312 358 402 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 478 312 583 402 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 699 312 804 402 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel metal1 969 196 1036 678 0 FreeSans 200 0 0 0 Y
port 9 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
