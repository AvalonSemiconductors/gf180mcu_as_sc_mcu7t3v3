magic
tech gf180mcuD
magscale 1 10
timestamp 1751882821
<< nwell >>
rect -86 354 1542 870
<< pwell >>
rect -86 -86 1542 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
<< ndiff >>
rect 28 255 116 268
rect 28 81 41 255
rect 87 81 116 255
rect 28 68 116 81
rect 172 242 276 268
rect 172 196 201 242
rect 247 196 276 242
rect 172 68 276 196
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 242 596 268
rect 492 196 521 242
rect 567 196 596 242
rect 492 68 596 196
rect 652 127 756 268
rect 652 81 681 127
rect 727 81 756 127
rect 652 68 756 81
rect 812 242 916 268
rect 812 196 841 242
rect 887 196 916 242
rect 812 68 916 196
rect 972 127 1076 268
rect 972 81 1001 127
rect 1047 81 1076 127
rect 972 68 1076 81
rect 1132 242 1236 268
rect 1132 196 1161 242
rect 1207 196 1236 242
rect 1132 68 1236 196
rect 1292 255 1428 268
rect 1292 81 1321 255
rect 1367 81 1428 255
rect 1292 68 1428 81
<< pdiff >>
rect 28 667 116 716
rect 28 480 41 667
rect 87 480 116 667
rect 28 440 116 480
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 526 436 716
rect 332 480 361 526
rect 407 480 436 526
rect 332 440 436 480
rect 492 703 596 716
rect 492 657 521 703
rect 567 657 596 703
rect 492 440 596 657
rect 652 667 756 716
rect 652 480 681 667
rect 727 480 756 667
rect 652 440 756 480
rect 812 550 916 716
rect 812 504 841 550
rect 887 504 916 550
rect 812 440 916 504
rect 972 678 1076 716
rect 972 632 1001 678
rect 1047 632 1076 678
rect 972 440 1076 632
rect 1132 550 1236 716
rect 1132 504 1161 550
rect 1207 504 1236 550
rect 1132 440 1236 504
rect 1292 678 1428 716
rect 1292 632 1321 678
rect 1367 632 1428 678
rect 1292 440 1428 632
<< ndiffc >>
rect 41 81 87 255
rect 201 196 247 242
rect 361 81 407 127
rect 521 196 567 242
rect 681 81 727 127
rect 841 196 887 242
rect 1001 81 1047 127
rect 1161 196 1207 242
rect 1321 81 1367 255
<< pdiffc >>
rect 41 480 87 667
rect 201 657 247 703
rect 361 480 407 526
rect 521 657 567 703
rect 681 480 727 667
rect 841 504 887 550
rect 1001 632 1047 678
rect 1161 504 1207 550
rect 1321 632 1367 678
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 116 393 172 440
rect 276 393 332 440
rect 436 393 492 440
rect 596 393 652 440
rect 116 379 652 393
rect 116 333 129 379
rect 639 333 652 379
rect 116 317 652 333
rect 116 268 172 317
rect 276 268 332 317
rect 436 268 492 317
rect 596 268 652 317
rect 756 393 812 440
rect 916 393 972 440
rect 1076 393 1132 440
rect 1236 393 1292 440
rect 756 379 1294 393
rect 756 333 771 379
rect 1095 333 1294 379
rect 756 317 1294 333
rect 756 268 812 317
rect 916 268 972 317
rect 1076 268 1132 317
rect 1236 268 1292 317
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
<< polycontact >>
rect 129 333 639 379
rect 771 333 1095 379
<< metal1 >>
rect 0 724 1456 844
rect 201 703 247 724
rect 41 667 87 678
rect 201 646 247 657
rect 521 703 567 724
rect 521 646 567 657
rect 681 667 1001 678
rect 87 480 361 526
rect 407 480 681 526
rect 727 632 1001 667
rect 1047 632 1321 678
rect 1367 632 1378 678
rect 1141 550 1227 553
rect 727 480 738 526
rect 795 504 841 550
rect 887 504 1161 550
rect 1207 504 1227 550
rect 41 464 87 480
rect 116 379 652 399
rect 116 333 129 379
rect 639 333 652 379
rect 116 313 652 333
rect 771 379 1095 397
rect 771 313 1095 333
rect 41 255 87 274
rect 1141 242 1227 504
rect 146 196 201 242
rect 247 196 521 242
rect 567 196 841 242
rect 887 196 1161 242
rect 1207 196 1227 242
rect 1321 255 1367 274
rect 41 60 87 81
rect 361 127 407 138
rect 361 60 407 81
rect 681 127 727 138
rect 681 60 727 81
rect 1001 127 1047 138
rect 1001 60 1047 81
rect 1321 60 1367 81
rect 0 -60 1456 60
<< labels >>
flabel metal1 s 0 724 1456 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1456 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 1141 196 1227 553 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 116 313 652 399 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 771 313 1095 397 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1472 354
string MASKHINTS_PPLUS -16 354 1472 830
<< end >>
