VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_12
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 0.205 2.850 0.435 3.620 ;
        RECT 1.805 2.765 2.035 3.620 ;
        RECT 3.405 2.770 3.635 3.620 ;
        RECT 5.005 2.770 5.235 3.620 ;
        RECT 6.605 2.765 6.835 3.620 ;
        RECT 8.205 2.265 8.435 3.620 ;
        RECT 9.820 2.265 10.050 3.620 ;
        RECT 11.420 2.265 11.650 3.620 ;
        RECT 13.020 2.265 13.250 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.840 ;
        RECT 1.805 0.300 2.035 0.710 ;
        RECT 3.405 0.300 3.635 0.710 ;
        RECT 5.005 0.300 5.235 0.710 ;
        RECT 6.605 0.300 6.835 0.710 ;
        RECT 8.205 0.300 8.435 1.300 ;
        RECT 9.820 0.300 10.050 1.300 ;
        RECT 11.420 0.300 11.650 1.300 ;
        RECT 13.020 0.300 13.250 1.300 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 1.570 3.145 2.075 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.461300 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 2.535 4.435 3.390 ;
        RECT 5.805 2.535 6.035 3.390 ;
        RECT 7.405 2.535 7.635 3.390 ;
        RECT 4.205 2.305 7.635 2.535 ;
        RECT 7.405 2.035 7.635 2.305 ;
        RECT 9.020 2.035 9.250 3.390 ;
        RECT 10.620 2.035 10.850 3.390 ;
        RECT 12.220 2.035 12.450 3.390 ;
        RECT 7.405 1.530 12.450 2.035 ;
        RECT 7.405 1.330 7.635 1.530 ;
        RECT 4.205 1.100 7.635 1.330 ;
        RECT 4.205 0.990 4.435 1.100 ;
        RECT 5.805 0.990 6.035 1.100 ;
        RECT 7.405 0.990 7.635 1.100 ;
        RECT 9.020 0.990 9.250 1.530 ;
        RECT 10.620 0.990 10.850 1.530 ;
        RECT 12.220 0.990 12.450 1.530 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.535 1.235 3.390 ;
        RECT 2.605 2.535 2.835 3.390 ;
        RECT 1.005 2.305 3.605 2.535 ;
        RECT 3.375 1.920 3.605 2.305 ;
        RECT 3.375 1.630 7.175 1.920 ;
        RECT 3.375 1.330 3.605 1.630 ;
        RECT 1.005 1.100 3.605 1.330 ;
        RECT 1.005 0.990 1.235 1.100 ;
        RECT 2.605 0.990 2.835 1.100 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_12


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.660 2.265 2.890 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.660 0.300 2.890 1.400 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.570 0.675 2.285 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.530 2.200 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.895 0.435 3.380 ;
        RECT 0.205 2.665 1.330 2.895 ;
        RECT 1.100 2.030 1.330 2.665 ;
        RECT 1.100 1.575 1.395 2.030 ;
        RECT 1.100 1.175 1.330 1.575 ;
        RECT 0.205 0.945 1.330 1.175 ;
        RECT 0.205 0.795 0.435 0.945 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.205 2.140 4.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 4.205 0.300 4.435 1.370 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.570 0.675 2.285 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 2.040 2.200 3.390 ;
        RECT 3.405 2.040 3.800 3.390 ;
        RECT 1.805 1.755 3.800 2.040 ;
        RECT 1.805 0.530 2.200 1.755 ;
        RECT 3.405 0.530 3.800 1.755 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.895 0.435 3.380 ;
        RECT 0.205 2.665 1.330 2.895 ;
        RECT 1.100 2.030 1.330 2.665 ;
        RECT 1.100 1.575 1.395 2.030 ;
        RECT 1.100 1.175 1.330 1.575 ;
        RECT 0.205 0.945 1.330 1.175 ;
        RECT 0.205 0.795 0.435 0.945 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_8
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.205 3.185 0.435 3.620 ;
        RECT 1.805 2.265 2.035 3.620 ;
        RECT 3.405 2.180 3.635 3.620 ;
        RECT 5.005 2.210 5.235 3.620 ;
        RECT 6.605 2.210 6.835 3.620 ;
        RECT 8.205 2.210 8.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.735 ;
        RECT 1.805 0.300 2.035 1.275 ;
        RECT 3.405 0.300 3.635 1.370 ;
        RECT 5.005 0.300 5.235 1.340 ;
        RECT 6.605 0.300 6.835 1.340 ;
        RECT 8.205 0.300 8.435 1.325 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 2.060 0.585 2.405 ;
        RECT 0.205 1.610 0.770 2.060 ;
        RECT 0.205 1.455 0.585 1.610 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.283200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 1.980 4.435 3.390 ;
        RECT 5.805 1.980 6.035 3.390 ;
        RECT 7.405 1.980 7.635 3.390 ;
        RECT 9.005 1.980 9.235 3.390 ;
        RECT 4.205 1.570 9.235 1.980 ;
        RECT 4.205 0.990 4.435 1.570 ;
        RECT 5.805 0.990 6.035 1.570 ;
        RECT 7.405 0.990 7.635 1.570 ;
        RECT 9.005 0.990 9.235 1.570 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.035 1.235 3.390 ;
        RECT 2.605 2.035 2.835 3.390 ;
        RECT 1.005 1.995 2.835 2.035 ;
        RECT 1.005 1.935 3.065 1.995 ;
        RECT 1.005 1.805 3.975 1.935 ;
        RECT 1.005 0.990 1.235 1.805 ;
        RECT 2.605 1.660 3.975 1.805 ;
        RECT 2.605 1.610 3.065 1.660 ;
        RECT 2.605 0.990 2.835 1.610 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__clkbuff_12
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__clkbuff_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 0.205 2.850 0.435 3.620 ;
        RECT 1.805 2.765 2.035 3.620 ;
        RECT 3.405 2.770 3.635 3.620 ;
        RECT 5.005 2.770 5.235 3.620 ;
        RECT 6.605 2.765 6.835 3.620 ;
        RECT 8.205 2.265 8.435 3.620 ;
        RECT 9.820 2.265 10.050 3.620 ;
        RECT 11.420 2.265 11.650 3.620 ;
        RECT 13.020 2.265 13.250 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.700 ;
        RECT 1.805 0.300 2.035 0.710 ;
        RECT 3.405 0.300 3.635 0.710 ;
        RECT 5.005 0.300 5.235 0.710 ;
        RECT 6.605 0.300 6.835 0.710 ;
        RECT 8.205 0.300 8.435 0.690 ;
        RECT 9.820 0.300 10.050 0.690 ;
        RECT 11.420 0.300 11.650 0.690 ;
        RECT 13.020 0.300 13.250 0.690 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 1.570 3.145 2.075 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 2.535 4.435 3.390 ;
        RECT 5.805 2.535 6.035 3.390 ;
        RECT 7.405 2.535 7.635 3.390 ;
        RECT 4.205 2.305 7.635 2.535 ;
        RECT 7.405 2.035 7.635 2.305 ;
        RECT 9.020 2.035 9.250 3.390 ;
        RECT 10.620 2.035 10.850 3.390 ;
        RECT 12.220 2.035 12.450 3.390 ;
        RECT 7.405 1.530 12.450 2.035 ;
        RECT 7.405 1.330 7.635 1.530 ;
        RECT 4.205 1.100 7.635 1.330 ;
        RECT 4.205 0.530 4.435 1.100 ;
        RECT 5.805 0.530 6.035 1.100 ;
        RECT 7.405 0.530 7.635 1.100 ;
        RECT 9.020 0.530 9.250 1.530 ;
        RECT 10.620 0.530 10.850 1.530 ;
        RECT 12.220 0.530 12.450 1.530 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.535 1.235 3.390 ;
        RECT 2.605 2.535 2.835 3.390 ;
        RECT 1.005 2.305 3.605 2.535 ;
        RECT 3.375 1.920 3.605 2.305 ;
        RECT 3.375 1.630 7.175 1.920 ;
        RECT 3.375 1.330 3.605 1.630 ;
        RECT 1.005 1.100 3.605 1.330 ;
        RECT 1.005 0.530 1.235 1.100 ;
        RECT 2.605 0.530 2.835 1.100 ;
  END
END gf180mcu_as_sc_mcu7t3v3__clkbuff_12


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__clkbuff_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__clkbuff_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.205 2.140 4.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 4.205 0.300 4.435 0.730 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.570 0.675 2.285 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.184000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 2.040 2.200 3.390 ;
        RECT 3.405 2.040 3.800 3.390 ;
        RECT 1.805 1.755 3.800 2.040 ;
        RECT 1.805 0.530 2.200 1.755 ;
        RECT 3.405 0.530 3.800 1.755 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.895 0.435 3.380 ;
        RECT 0.205 2.665 1.330 2.895 ;
        RECT 1.100 2.030 1.330 2.665 ;
        RECT 1.100 1.575 1.395 2.030 ;
        RECT 1.100 1.175 1.330 1.575 ;
        RECT 0.205 0.945 1.330 1.175 ;
        RECT 0.205 0.530 0.435 0.945 ;
  END
END gf180mcu_as_sc_mcu7t3v3__clkbuff_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__clkbuff_8
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__clkbuff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.205 3.185 0.435 3.620 ;
        RECT 1.805 2.265 2.035 3.620 ;
        RECT 3.405 2.180 3.635 3.620 ;
        RECT 5.005 2.210 5.235 3.620 ;
        RECT 6.605 2.210 6.835 3.620 ;
        RECT 8.205 2.210 8.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.735 ;
        RECT 1.805 0.300 2.035 0.700 ;
        RECT 3.405 0.300 3.635 0.795 ;
        RECT 5.005 0.300 5.235 0.765 ;
        RECT 6.605 0.300 6.835 0.765 ;
        RECT 8.205 0.300 8.435 0.750 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.764000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 2.060 0.585 2.405 ;
        RECT 0.205 1.610 0.770 2.060 ;
        RECT 0.205 1.455 0.585 1.610 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.544000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 1.980 4.435 3.390 ;
        RECT 5.805 1.980 6.035 3.390 ;
        RECT 7.405 1.980 7.635 3.390 ;
        RECT 9.005 1.980 9.235 3.390 ;
        RECT 4.205 1.570 9.235 1.980 ;
        RECT 4.205 0.710 4.435 1.570 ;
        RECT 5.805 0.710 6.035 1.570 ;
        RECT 7.405 0.710 7.635 1.570 ;
        RECT 9.005 0.710 9.235 1.570 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.035 1.235 3.390 ;
        RECT 2.605 2.035 2.835 3.390 ;
        RECT 1.005 1.995 2.835 2.035 ;
        RECT 1.005 1.935 3.065 1.995 ;
        RECT 1.005 1.805 3.975 1.935 ;
        RECT 1.005 0.710 1.235 1.805 ;
        RECT 2.605 1.660 3.975 1.805 ;
        RECT 2.605 1.610 3.065 1.660 ;
        RECT 2.605 0.710 2.835 1.610 ;
  END
END gf180mcu_as_sc_mcu7t3v3__clkbuff_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__decap_16
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__decap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 8.525 2.555 8.755 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.740 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.240 1.735 0.470 3.390 ;
        RECT 8.020 2.095 8.755 2.325 ;
        RECT 0.240 1.500 1.040 1.735 ;
        RECT 0.650 1.440 1.040 1.500 ;
        RECT 8.525 0.980 8.755 2.095 ;
  END
END gf180mcu_as_sc_mcu7t3v3__decap_16


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__decap_4
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 1.805 2.565 2.035 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.740 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.240 1.735 0.470 3.390 ;
        RECT 1.305 2.090 2.035 2.335 ;
        RECT 0.240 1.500 1.040 1.735 ;
        RECT 0.650 1.440 1.040 1.500 ;
        RECT 1.805 0.530 2.035 2.090 ;
  END
END gf180mcu_as_sc_mcu7t3v3__decap_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__decap_8
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__decap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 4.045 2.565 4.275 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.740 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.240 1.735 0.470 3.390 ;
        RECT 3.520 2.095 4.275 2.335 ;
        RECT 0.240 1.500 1.040 1.735 ;
        RECT 0.650 1.440 1.040 1.500 ;
        RECT 4.045 0.980 4.275 2.095 ;
  END
END gf180mcu_as_sc_mcu7t3v3__decap_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__dfxtp_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.490 3.230 2.720 3.620 ;
        RECT 7.000 3.230 7.230 3.620 ;
        RECT 11.360 3.230 11.590 3.620 ;
        RECT 12.910 2.145 13.140 3.620 ;
        RECT 14.510 2.145 14.740 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 15.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.490 0.300 2.720 0.690 ;
        RECT 7.000 0.300 7.230 0.690 ;
        RECT 11.360 0.300 11.590 0.690 ;
        RECT 12.910 0.300 13.140 1.390 ;
        RECT 14.510 0.300 14.740 1.385 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 1.600 0.860 2.060 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.985 1.630 4.430 2.930 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.615 0.990 14.045 2.550 ;
    END
  END Q
  OBS
      LAYER Metal1 ;
        RECT 2.970 3.160 6.205 3.390 ;
        RECT 2.970 3.000 3.200 3.160 ;
        RECT 0.205 2.935 0.445 2.995 ;
        RECT 1.105 2.935 3.200 3.000 ;
        RECT 0.205 2.770 3.200 2.935 ;
        RECT 0.205 2.705 1.335 2.770 ;
        RECT 0.205 2.650 0.445 2.705 ;
        RECT 1.105 1.985 1.335 2.705 ;
        RECT 1.745 2.265 2.095 2.495 ;
        RECT 1.805 2.000 2.035 2.265 ;
        RECT 1.105 1.605 1.405 1.985 ;
        RECT 1.805 1.770 3.680 2.000 ;
        RECT 0.205 1.275 0.435 1.330 ;
        RECT 1.105 1.275 1.335 1.605 ;
        RECT 0.205 1.045 1.335 1.275 ;
        RECT 0.205 0.990 0.435 1.045 ;
        RECT 1.805 0.990 2.035 1.770 ;
        RECT 3.375 1.640 3.680 1.770 ;
        RECT 3.450 0.760 3.680 1.640 ;
        RECT 4.660 1.400 4.890 2.550 ;
        RECT 5.120 1.630 5.350 3.160 ;
        RECT 5.925 3.090 6.205 3.160 ;
        RECT 5.925 2.755 6.305 3.090 ;
        RECT 8.320 3.005 10.620 3.235 ;
        RECT 5.580 2.295 7.530 2.525 ;
        RECT 5.580 1.400 5.810 2.295 ;
        RECT 6.045 1.990 6.325 2.025 ;
        RECT 4.660 1.170 5.810 1.400 ;
        RECT 6.040 1.645 6.325 1.990 ;
        RECT 4.660 0.990 4.890 1.170 ;
        RECT 6.040 0.760 6.270 1.645 ;
        RECT 6.625 1.640 6.885 1.990 ;
        RECT 6.655 1.220 6.885 1.640 ;
        RECT 7.300 1.625 7.530 2.295 ;
        RECT 7.800 1.220 8.030 2.550 ;
        RECT 8.320 1.985 8.550 3.005 ;
        RECT 8.260 1.595 8.640 1.985 ;
        RECT 8.870 1.560 9.190 2.025 ;
        RECT 6.655 0.990 8.030 1.220 ;
        RECT 9.420 1.150 9.650 2.550 ;
        RECT 10.390 1.625 10.620 3.005 ;
        RECT 12.270 2.500 12.500 3.390 ;
        RECT 11.010 2.270 12.500 2.500 ;
        RECT 11.010 1.625 11.240 2.270 ;
        RECT 12.270 1.980 12.500 2.270 ;
        RECT 11.810 1.150 12.040 1.980 ;
        RECT 9.420 0.920 12.040 1.150 ;
        RECT 12.270 1.620 12.650 1.980 ;
        RECT 12.270 0.990 12.500 1.620 ;
        RECT 3.450 0.530 6.270 0.760 ;
      LAYER Metal2 ;
        RECT 5.915 2.760 9.200 3.040 ;
        RECT 6.045 1.975 6.325 2.025 ;
        RECT 6.035 1.695 8.640 1.975 ;
        RECT 6.045 1.645 6.325 1.695 ;
        RECT 8.920 1.640 9.200 2.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__dfxtp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 1.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.330 0.805 0.630 2.750 ;
    END
  END DIODE
END gf180mcu_as_sc_mcu7t3v3__diode_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_1
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 0.560 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 0.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 0.990 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 0.560 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_1


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_2
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 1.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_4
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_8
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__inv_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.205 2.355 0.435 3.620 ;
        RECT 1.805 2.295 2.035 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.235 ;
        RECT 1.805 0.300 2.035 1.235 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.255 1.235 3.385 ;
        RECT 1.005 1.260 1.350 2.255 ;
        RECT 1.005 0.530 1.235 1.260 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.590 0.775 2.125 ;
    END
  END A
END gf180mcu_as_sc_mcu7t3v3__inv_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__inv_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 0.205 2.355 0.435 3.620 ;
        RECT 1.805 2.295 2.035 3.620 ;
        RECT 3.405 2.175 3.635 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.235 ;
        RECT 1.805 0.300 2.035 1.235 ;
        RECT 3.405 0.300 3.635 1.395 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.255 1.235 3.385 ;
        RECT 1.005 1.935 1.350 2.255 ;
        RECT 2.605 1.935 2.835 3.385 ;
        RECT 1.005 1.705 2.835 1.935 ;
        RECT 1.005 1.260 1.350 1.705 ;
        RECT 1.005 0.990 1.235 1.260 ;
        RECT 2.605 0.990 2.835 1.705 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.590 0.775 2.125 ;
    END
  END A
END gf180mcu_as_sc_mcu7t3v3__inv_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 0.205 2.840 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.410 3.230 3.640 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.955200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 3.000 1.235 3.160 ;
        RECT 2.605 3.000 2.835 3.160 ;
        RECT 1.005 2.770 3.635 3.000 ;
        RECT 2.605 1.320 2.835 1.330 ;
        RECT 3.165 1.320 3.635 2.770 ;
        RECT 2.605 1.050 3.635 1.320 ;
        RECT 2.605 0.990 2.835 1.050 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.130 1.610 2.935 2.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 1.615 1.660 2.020 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 0.205 0.920 2.035 1.150 ;
        RECT 0.205 0.805 0.435 0.920 ;
        RECT 1.805 0.760 2.035 0.920 ;
        RECT 1.805 0.530 3.690 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nor2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.757600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.545 2.285 3.635 2.555 ;
        RECT 2.605 1.320 2.835 1.330 ;
        RECT 3.165 1.320 3.635 2.285 ;
        RECT 2.605 1.275 3.635 1.320 ;
        RECT 1.005 1.050 3.635 1.275 ;
        RECT 1.005 1.045 2.835 1.050 ;
        RECT 1.005 0.935 1.235 1.045 ;
        RECT 2.605 0.990 2.835 1.045 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.130 1.610 2.935 2.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 1.615 1.660 2.020 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.750 3.160 3.690 3.390 ;
        RECT 0.205 2.925 0.435 3.040 ;
        RECT 1.750 2.925 1.980 3.160 ;
        RECT 0.205 2.695 1.980 2.925 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nor2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__tap_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 1.550 4.350 ;
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
        RECT 0.375 1.930 0.715 3.620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.770 ;
      LAYER Metal1 ;
        RECT 0.375 0.300 0.715 1.510 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__tap_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__tieh_4
  CLASS CORE TIEHIGH ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__tieh_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.205 2.220 0.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.375 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN ONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.190 1.365 3.390 ;
    END
  END ONE
  OBS
      LAYER Metal1 ;
        RECT 0.570 1.660 1.235 1.895 ;
        RECT 1.005 0.530 1.235 1.660 ;
  END
END gf180mcu_as_sc_mcu7t3v3__tieh_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__tiel_4
  CLASS CORE TIELOW ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__tiel_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.205 2.220 0.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.375 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN ZERO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.920 0.530 1.280 1.425 ;
    END
  END ZERO
  OBS
      LAYER Metal1 ;
        RECT 1.005 1.895 1.235 3.390 ;
        RECT 0.570 1.660 1.235 1.895 ;
  END
END gf180mcu_as_sc_mcu7t3v3__tiel_4


END LIBRARY
