magic
tech gf180mcuD
magscale 1 10
timestamp 1751740063
<< nwell >>
rect -86 354 870 870
<< pwell >>
rect -86 -86 870 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 244 276 268
rect 172 198 201 244
rect 247 198 276 244
rect 172 68 276 198
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 255 596 268
rect 492 209 521 255
rect 567 209 596 255
rect 492 68 596 209
rect 652 127 755 268
rect 652 81 681 127
rect 727 81 755 127
rect 652 68 755 81
<< pdiff >>
rect 28 597 116 716
rect 28 551 41 597
rect 87 551 116 597
rect 28 440 116 551
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 678 436 716
rect 332 632 361 678
rect 407 632 436 678
rect 332 440 436 632
rect 492 503 596 716
rect 492 457 521 503
rect 567 457 596 503
rect 492 440 596 457
rect 652 678 756 716
rect 652 632 681 678
rect 727 632 756 678
rect 652 440 756 632
<< ndiffc >>
rect 41 81 87 127
rect 201 198 247 244
rect 361 81 407 127
rect 521 209 567 255
rect 681 81 727 127
<< pdiffc >>
rect 41 551 87 597
rect 201 657 247 703
rect 361 632 407 678
rect 521 457 567 503
rect 681 632 727 678
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 116 404 172 440
rect 276 404 332 440
rect 100 388 332 404
rect 436 403 492 440
rect 596 403 652 440
rect 100 342 114 388
rect 319 342 332 388
rect 100 323 332 342
rect 116 268 172 323
rect 276 268 332 323
rect 426 387 652 403
rect 426 341 439 387
rect 587 341 652 387
rect 426 322 652 341
rect 436 268 492 322
rect 596 268 652 322
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
<< polycontact >>
rect 114 342 319 388
rect 439 341 587 387
<< metal1 >>
rect 0 724 784 844
rect 201 703 247 724
rect 201 646 247 657
rect 350 632 361 678
rect 407 632 681 678
rect 727 632 738 678
rect 41 597 87 608
rect 350 585 396 632
rect 87 551 396 585
rect 41 539 396 551
rect 509 503 727 511
rect 509 457 521 503
rect 567 457 727 503
rect 100 388 332 404
rect 100 342 114 388
rect 319 342 332 388
rect 100 323 332 342
rect 426 387 587 403
rect 426 341 439 387
rect 426 322 587 341
rect 521 264 567 266
rect 633 264 727 457
rect 521 255 727 264
rect 201 244 521 255
rect 247 209 521 244
rect 567 210 727 255
rect 521 198 567 209
rect 201 187 247 198
rect 41 127 87 138
rect 41 60 87 81
rect 361 127 407 138
rect 361 60 407 81
rect 681 127 727 138
rect 681 60 727 81
rect 0 -60 784 60
<< labels >>
flabel metal1 s 0 724 784 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 784 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 633 210 727 511 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 426 322 587 403 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 100 323 332 404 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 784 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 870 354
string MASKHINTS_PPLUS -86 354 870 870
<< end >>
