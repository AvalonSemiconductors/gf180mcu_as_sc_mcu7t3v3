VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__and2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 0.205 3.230 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 2.150 3.635 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 1.450 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.555 1.660 2.540 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.560 0.860 1.985 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.605 0.920 3.035 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.950 2.770 2.120 3.000 ;
        RECT 1.890 1.980 2.120 2.770 ;
        RECT 1.890 1.555 2.195 1.980 ;
        RECT 0.205 1.150 0.435 1.240 ;
        RECT 1.890 1.150 2.120 1.555 ;
        RECT 0.205 0.920 2.120 1.150 ;
        RECT 0.205 0.860 0.435 0.920 ;
  END
END gf180mcu_as_sc_mcu7t3v3__and2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__and2_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.205 3.230 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 2.150 3.635 3.620 ;
        RECT 5.005 2.150 5.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 1.450 ;
        RECT 5.005 0.300 5.235 1.450 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.555 1.660 2.540 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.560 0.860 1.985 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.605 1.920 2.835 3.390 ;
        RECT 4.205 1.920 4.600 3.390 ;
        RECT 2.605 1.690 4.600 1.920 ;
        RECT 2.605 0.920 2.835 1.690 ;
        RECT 4.205 0.920 4.600 1.690 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.950 2.770 2.120 3.000 ;
        RECT 1.890 1.980 2.120 2.770 ;
        RECT 1.890 1.555 2.195 1.980 ;
        RECT 0.205 1.150 0.435 1.240 ;
        RECT 1.890 1.150 2.120 1.555 ;
        RECT 0.205 0.920 2.120 1.150 ;
        RECT 0.205 0.860 0.435 0.920 ;
  END
END gf180mcu_as_sc_mcu7t3v3__and2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao211_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 1.005 3.190 1.235 3.620 ;
        RECT 4.045 2.260 4.275 3.620 ;
        RECT 5.645 2.460 5.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.730 ;
        RECT 2.605 0.300 2.835 0.730 ;
        RECT 4.045 0.300 4.275 0.730 ;
        RECT 5.645 0.300 5.875 0.730 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.330 1.550 0.715 2.265 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 1.320 1.615 2.255 ;
        RECT 1.230 0.595 1.575 1.320 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.030 1.570 2.415 2.260 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.830 1.535 3.215 2.290 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.815 0.840 5.125 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.960 0.435 3.175 ;
        RECT 1.805 2.960 2.035 3.160 ;
        RECT 0.205 2.730 2.035 2.960 ;
        RECT 3.405 2.750 3.635 3.390 ;
        RECT 3.405 2.520 3.700 2.750 ;
        RECT 3.470 1.955 3.700 2.520 ;
        RECT 3.470 1.575 4.440 1.955 ;
        RECT 3.470 1.190 3.700 1.575 ;
        RECT 1.805 0.960 3.700 1.190 ;
        RECT 1.805 0.735 2.035 0.960 ;
        RECT 3.405 0.790 3.700 0.960 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao211_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao211_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 1.005 3.190 1.235 3.620 ;
        RECT 4.045 2.260 4.275 3.620 ;
        RECT 5.645 2.260 5.875 3.620 ;
        RECT 7.245 2.260 7.475 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.730 ;
        RECT 2.605 0.300 2.835 0.730 ;
        RECT 4.045 0.300 4.275 0.730 ;
        RECT 5.645 0.300 5.875 0.730 ;
        RECT 7.245 0.300 7.475 0.730 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.330 1.550 0.715 2.265 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.230 1.320 1.615 2.255 ;
        RECT 1.230 0.595 1.575 1.320 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.030 1.570 2.415 2.260 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.830 1.535 3.215 2.290 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.815 1.935 5.125 3.390 ;
        RECT 6.415 1.935 6.725 3.390 ;
        RECT 4.815 1.600 6.725 1.935 ;
        RECT 4.815 0.840 5.125 1.600 ;
        RECT 6.415 0.840 6.725 1.600 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.960 0.435 3.175 ;
        RECT 1.805 2.960 2.035 3.160 ;
        RECT 0.205 2.730 2.035 2.960 ;
        RECT 3.405 2.750 3.635 3.390 ;
        RECT 3.405 2.520 3.700 2.750 ;
        RECT 3.470 1.955 3.700 2.520 ;
        RECT 3.470 1.575 4.440 1.955 ;
        RECT 3.470 1.190 3.700 1.575 ;
        RECT 1.805 0.960 3.700 1.190 ;
        RECT 1.805 0.735 2.035 0.960 ;
        RECT 3.405 0.790 3.700 0.960 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao211_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao21_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 3.245 2.145 3.475 3.620 ;
        RECT 4.930 2.145 5.160 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 2.605 0.300 3.475 0.690 ;
        RECT 4.930 0.300 5.160 1.380 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.439900 ;
    PORT
      LAYER Metal1 ;
        RECT 4.130 0.990 4.450 3.380 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 1.580 0.860 2.360 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 1.580 1.660 1.965 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 1.580 2.460 1.965 ;
    END
  END C
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.975 0.435 3.100 ;
        RECT 1.805 2.975 2.035 3.045 ;
        RECT 0.205 2.745 2.035 2.975 ;
        RECT 0.205 2.665 0.435 2.745 ;
        RECT 1.805 2.670 2.035 2.745 ;
        RECT 2.605 2.475 2.835 3.390 ;
        RECT 2.605 2.225 2.925 2.475 ;
        RECT 2.695 1.885 2.925 2.225 ;
        RECT 2.695 1.655 3.900 1.885 ;
        RECT 2.695 1.240 2.925 1.655 ;
        RECT 1.745 1.010 2.925 1.240 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao21_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao21_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 3.245 2.145 3.475 3.620 ;
        RECT 4.930 2.145 5.160 3.620 ;
        RECT 6.530 2.145 6.760 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 2.605 0.300 3.475 0.690 ;
        RECT 4.930 0.300 5.160 1.380 ;
        RECT 6.530 0.300 6.760 1.380 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.677500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.130 1.890 4.450 3.380 ;
        RECT 5.730 1.890 6.050 3.380 ;
        RECT 4.130 1.660 6.050 1.890 ;
        RECT 4.130 0.990 4.450 1.660 ;
        RECT 5.730 0.990 6.050 1.660 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 1.580 0.860 2.360 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.200 1.580 1.660 1.965 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.000 1.580 2.460 1.965 ;
    END
  END C
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.975 0.435 3.100 ;
        RECT 1.805 2.975 2.035 3.045 ;
        RECT 0.205 2.745 2.035 2.975 ;
        RECT 0.205 2.665 0.435 2.745 ;
        RECT 1.805 2.670 2.035 2.745 ;
        RECT 2.605 2.475 2.835 3.390 ;
        RECT 2.605 2.225 2.925 2.475 ;
        RECT 2.695 1.885 2.925 2.225 ;
        RECT 2.695 1.655 3.900 1.885 ;
        RECT 2.695 1.240 2.925 1.655 ;
        RECT 1.745 1.010 2.925 1.240 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao21_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao21b_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao21b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
        RECT 0.425 2.515 0.655 3.620 ;
        RECT 2.685 3.230 2.915 3.620 ;
        RECT 4.285 3.230 4.515 3.620 ;
        RECT 7.325 3.230 7.555 3.620 ;
        RECT 8.925 3.230 9.155 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 9.950 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.950 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 0.300 0.645 0.690 ;
        RECT 1.885 0.300 2.115 0.690 ;
        RECT 5.085 0.300 5.315 0.690 ;
        RECT 6.685 0.300 7.550 0.690 ;
        RECT 8.925 0.300 9.155 0.690 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 8.110 0.990 8.375 3.390 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.415 1.565 6.805 2.310 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 1.590 4.140 1.950 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.480 1.015 2.285 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.945 1.475 3.390 ;
        RECT 5.085 3.160 6.915 3.390 ;
        RECT 1.885 3.000 2.115 3.080 ;
        RECT 5.085 3.000 5.315 3.160 ;
        RECT 1.885 2.770 5.315 3.000 ;
        RECT 6.685 2.970 6.915 3.160 ;
        RECT 1.885 2.695 2.115 2.770 ;
        RECT 2.325 2.310 4.770 2.540 ;
        RECT 2.325 1.955 2.555 2.310 ;
        RECT 2.135 1.945 2.555 1.955 ;
        RECT 1.245 1.595 2.555 1.945 ;
        RECT 1.245 0.985 1.475 1.595 ;
        RECT 2.135 1.590 2.555 1.595 ;
        RECT 4.540 1.930 4.770 2.310 ;
        RECT 4.540 1.570 4.945 1.930 ;
        RECT 5.825 1.255 6.115 2.620 ;
        RECT 7.485 1.545 7.870 1.945 ;
        RECT 7.485 1.255 7.715 1.545 ;
        RECT 3.360 1.025 7.715 1.255 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao21b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao21b_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao21b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.200 4.220 ;
        RECT 0.425 2.515 0.655 3.620 ;
        RECT 2.685 3.230 2.915 3.620 ;
        RECT 4.285 3.230 4.515 3.620 ;
        RECT 7.325 3.230 7.555 3.620 ;
        RECT 8.925 3.230 9.155 3.620 ;
        RECT 10.525 3.230 10.755 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 11.630 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.630 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 0.300 0.645 0.690 ;
        RECT 1.885 0.300 2.115 0.690 ;
        RECT 5.085 0.300 5.315 0.690 ;
        RECT 6.685 0.300 7.550 0.690 ;
        RECT 8.925 0.300 9.155 0.690 ;
        RECT 10.525 0.300 10.755 0.690 ;
        RECT 0.000 -0.300 11.200 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 8.110 1.895 8.375 3.390 ;
        RECT 9.700 1.895 9.965 3.390 ;
        RECT 8.110 1.645 9.965 1.895 ;
        RECT 8.110 0.990 8.375 1.645 ;
        RECT 9.700 0.990 9.965 1.645 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.415 1.565 6.805 2.310 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 1.590 4.140 1.950 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.480 1.015 2.285 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.945 1.475 3.390 ;
        RECT 5.085 3.160 6.915 3.390 ;
        RECT 1.885 3.000 2.115 3.080 ;
        RECT 5.085 3.000 5.315 3.160 ;
        RECT 1.885 2.770 5.315 3.000 ;
        RECT 6.685 2.970 6.915 3.160 ;
        RECT 1.885 2.695 2.115 2.770 ;
        RECT 2.325 2.310 4.770 2.540 ;
        RECT 2.325 1.955 2.555 2.310 ;
        RECT 2.135 1.945 2.555 1.955 ;
        RECT 1.245 1.595 2.555 1.945 ;
        RECT 1.245 0.985 1.475 1.595 ;
        RECT 2.135 1.590 2.555 1.595 ;
        RECT 4.540 1.930 4.770 2.310 ;
        RECT 4.540 1.570 4.945 1.930 ;
        RECT 5.825 1.255 6.115 2.620 ;
        RECT 7.485 1.545 7.870 1.945 ;
        RECT 7.485 1.255 7.715 1.545 ;
        RECT 3.360 1.025 7.715 1.255 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao21b_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao22_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 2.445 3.230 2.675 3.620 ;
        RECT 4.045 3.230 4.275 3.620 ;
        RECT 5.645 2.155 5.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 4.045 0.300 4.275 0.690 ;
        RECT 5.645 0.300 5.875 1.385 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.335 1.560 0.860 2.010 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.560 1.790 2.010 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.560 2.915 2.010 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.495 1.560 4.020 2.010 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.845 0.980 5.180 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.160 2.090 3.390 ;
        RECT 0.205 2.470 0.435 3.160 ;
        RECT 3.245 2.930 3.475 3.160 ;
        RECT 0.900 2.700 3.475 2.930 ;
        RECT 0.205 2.240 4.590 2.470 ;
        RECT 4.360 1.245 4.590 2.240 ;
        RECT 3.250 1.015 4.590 1.245 ;
        RECT 3.250 0.760 3.480 1.015 ;
        RECT 1.635 0.530 3.480 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao22_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao22_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 2.445 3.230 2.675 3.620 ;
        RECT 4.045 3.230 4.275 3.620 ;
        RECT 5.645 2.155 5.875 3.620 ;
        RECT 7.245 2.155 7.475 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 4.045 0.300 4.275 0.690 ;
        RECT 5.645 0.300 5.875 1.385 ;
        RECT 7.245 0.300 7.475 1.385 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.335 1.560 0.860 2.010 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.560 1.790 2.010 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.390 1.560 2.915 2.010 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.495 1.560 4.020 2.010 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.845 1.880 5.180 3.390 ;
        RECT 6.445 1.880 6.780 3.390 ;
        RECT 4.845 1.650 6.780 1.880 ;
        RECT 4.845 0.980 5.180 1.650 ;
        RECT 6.445 0.980 6.780 1.650 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.160 2.090 3.390 ;
        RECT 0.205 2.470 0.435 3.160 ;
        RECT 3.245 2.930 3.475 3.160 ;
        RECT 0.900 2.700 3.475 2.930 ;
        RECT 0.205 2.240 4.590 2.470 ;
        RECT 4.360 1.245 4.590 2.240 ;
        RECT 3.250 1.015 4.590 1.245 ;
        RECT 3.250 0.760 3.480 1.015 ;
        RECT 1.635 0.530 3.480 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao22_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao31_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 3.230 3.635 3.620 ;
        RECT 5.005 2.180 5.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 5.005 0.300 5.235 1.370 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 1.585 1.085 2.435 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.380 1.585 1.800 2.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.180 1.150 2.600 2.000 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.980 1.585 3.320 2.105 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 0.990 4.545 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 1.150 0.435 3.390 ;
        RECT 0.950 2.770 2.900 3.000 ;
        RECT 3.745 1.915 3.975 1.970 ;
        RECT 3.630 1.630 3.975 1.915 ;
        RECT 3.630 1.150 3.860 1.630 ;
        RECT 0.205 0.920 1.235 1.150 ;
        RECT 1.005 0.760 1.235 0.920 ;
        RECT 2.945 0.920 3.860 1.150 ;
        RECT 2.945 0.760 3.175 0.920 ;
        RECT 1.005 0.530 3.175 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao31_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__ao31_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__ao31_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 3.230 3.635 3.620 ;
        RECT 5.005 2.180 5.235 3.620 ;
        RECT 6.605 2.180 6.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 5.005 0.300 5.235 1.370 ;
        RECT 6.605 0.300 6.835 1.370 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 1.585 1.085 2.435 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.380 1.585 1.800 2.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.180 1.150 2.600 2.000 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 2.980 1.585 3.320 2.105 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 1.910 4.545 3.390 ;
        RECT 5.805 1.910 6.145 3.390 ;
        RECT 4.205 1.680 6.145 1.910 ;
        RECT 4.205 0.990 4.545 1.680 ;
        RECT 5.805 0.990 6.145 1.680 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 1.150 0.435 3.390 ;
        RECT 0.950 2.770 2.900 3.000 ;
        RECT 3.745 1.915 3.975 1.970 ;
        RECT 3.630 1.630 3.975 1.915 ;
        RECT 3.630 1.150 3.860 1.630 ;
        RECT 0.205 0.920 1.235 1.150 ;
        RECT 1.005 0.760 1.235 0.920 ;
        RECT 2.945 0.920 3.860 1.150 ;
        RECT 2.945 0.760 3.175 0.920 ;
        RECT 1.005 0.530 3.175 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__ao31_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi211_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.205 2.335 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 3.230 3.635 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 4.045 0.300 4.275 0.690 ;
        RECT 5.645 0.300 5.875 0.690 ;
        RECT 7.245 0.300 7.475 0.690 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 1.570 0.855 2.065 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.135 1.595 3.215 2.025 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.265 1.595 5.240 1.945 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.277600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.735 2.630 6.730 2.860 ;
        RECT 2.605 1.325 2.835 1.345 ;
        RECT 5.735 1.325 6.160 2.630 ;
        RECT 2.605 1.095 6.675 1.325 ;
        RECT 2.605 0.990 2.835 1.095 ;
        RECT 4.845 0.530 5.075 1.095 ;
        RECT 6.445 0.530 6.675 1.095 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.820 1.565 7.470 2.040 ;
    END
  END D
  OBS
      LAYER Metal1 ;
        RECT 3.990 3.160 7.530 3.390 ;
        RECT 2.605 2.685 5.130 2.850 ;
        RECT 0.950 2.620 5.130 2.685 ;
        RECT 0.950 2.455 2.835 2.620 ;
        RECT 0.205 0.965 2.035 1.195 ;
        RECT 0.205 0.775 0.435 0.965 ;
        RECT 1.805 0.760 2.035 0.965 ;
        RECT 1.805 0.530 3.690 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi211_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi211_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi211_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.205 3.230 4.435 3.620 ;
        RECT 5.805 3.230 6.035 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 6.605 0.300 6.835 0.690 ;
        RECT 8.205 0.300 8.435 0.690 ;
        RECT 9.805 0.300 10.035 0.690 ;
        RECT 11.405 0.300 11.635 0.690 ;
        RECT 13.005 0.300 13.235 0.690 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.125 2.215 6.435 2.445 ;
        RECT 2.125 1.975 2.460 2.215 ;
        RECT 0.580 1.575 2.460 1.975 ;
        RECT 6.205 1.570 6.435 2.215 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.980 1.565 5.565 1.960 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.980 1.565 8.885 1.955 ;
        RECT 12.485 1.590 12.900 1.940 ;
      LAYER Metal2 ;
        RECT 8.555 1.320 8.885 1.905 ;
        RECT 12.580 1.320 12.860 1.950 ;
        RECT 8.555 1.040 12.860 1.320 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 9.380 1.600 12.015 1.940 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.555200 ;
    PORT
      LAYER Metal1 ;
        RECT 9.750 2.745 12.370 2.975 ;
        RECT 12.140 2.700 12.370 2.745 ;
        RECT 12.140 2.470 13.475 2.700 ;
        RECT 13.130 1.220 13.475 2.470 ;
        RECT 3.350 0.990 13.475 1.220 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.000 0.435 3.390 ;
        RECT 6.605 3.160 8.595 3.390 ;
        RECT 6.605 3.000 6.835 3.160 ;
        RECT 0.205 2.770 6.835 3.000 ;
        RECT 8.205 2.955 8.595 3.160 ;
        RECT 12.915 2.930 13.235 3.390 ;
        RECT 7.350 2.470 7.690 2.495 ;
        RECT 10.550 2.470 10.890 2.495 ;
        RECT 7.350 2.240 10.890 2.470 ;
        RECT 1.005 0.920 2.835 1.150 ;
        RECT 1.005 0.790 1.235 0.920 ;
        RECT 2.605 0.760 2.835 0.920 ;
        RECT 2.605 0.530 6.095 0.760 ;
      LAYER Metal2 ;
        RECT 8.220 3.235 8.600 3.305 ;
        RECT 12.880 3.235 13.225 3.310 ;
        RECT 8.220 2.955 13.225 3.235 ;
        RECT 12.880 2.930 13.225 2.955 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi211_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi21_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi21_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 5.005 0.300 5.235 0.690 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.757600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.145 1.255 4.435 2.620 ;
        RECT 1.680 1.025 4.490 1.255 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.735 1.565 5.125 2.310 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.380 1.590 2.460 1.950 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 2.310 3.090 2.540 ;
        RECT 0.645 1.955 0.875 2.310 ;
        RECT 0.455 1.590 0.875 1.955 ;
        RECT 2.860 1.930 3.090 2.310 ;
        RECT 2.860 1.570 3.265 1.930 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 3.405 3.160 5.235 3.390 ;
        RECT 0.205 3.000 0.435 3.080 ;
        RECT 3.405 3.000 3.635 3.160 ;
        RECT 0.205 2.770 3.635 3.000 ;
        RECT 5.005 2.970 5.235 3.160 ;
        RECT 0.205 2.695 0.435 2.770 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi21_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi21_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi21_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.640 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.640 4.220 ;
        RECT 4.205 3.230 4.435 3.620 ;
        RECT 5.805 3.230 6.035 3.620 ;
        RECT 7.405 3.230 7.635 3.620 ;
        RECT 9.005 3.230 9.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 11.070 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 11.070 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 8.205 0.300 8.435 0.690 ;
        RECT 9.805 0.300 10.035 1.370 ;
        RECT 0.000 -0.300 10.640 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.515200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.935 2.265 3.095 2.495 ;
        RECT 2.750 1.275 3.095 2.265 ;
        RECT 0.805 1.045 6.895 1.275 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.380 1.590 2.520 1.955 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.760 2.310 8.010 2.540 ;
        RECT 3.760 1.955 3.990 2.310 ;
        RECT 3.565 1.590 3.990 1.955 ;
        RECT 7.780 1.955 8.010 2.310 ;
        RECT 7.780 1.590 9.660 1.955 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.580 1.590 7.260 1.955 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.105 3.690 3.335 ;
        RECT 0.205 2.870 0.435 3.105 ;
        RECT 3.460 3.000 3.690 3.105 ;
        RECT 9.805 3.000 10.035 3.300 ;
        RECT 3.460 2.770 10.035 3.000 ;
        RECT 7.405 0.990 9.235 1.220 ;
        RECT 7.405 0.760 7.635 0.990 ;
        RECT 4.100 0.530 7.635 0.760 ;
        RECT 9.005 0.655 9.235 0.990 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi21_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi21b_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi21b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 0.425 2.515 0.655 3.620 ;
        RECT 2.685 3.230 2.915 3.620 ;
        RECT 4.285 3.230 4.515 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 0.300 0.645 0.690 ;
        RECT 1.885 0.300 2.115 0.690 ;
        RECT 5.085 0.300 5.315 0.690 ;
        RECT 6.685 0.300 6.915 0.690 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.757600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.825 1.255 6.115 2.620 ;
        RECT 3.360 1.025 6.170 1.255 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.415 1.565 6.805 2.310 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.060 1.590 4.140 1.950 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 1.480 1.015 2.285 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.945 1.475 3.390 ;
        RECT 5.085 3.160 6.915 3.390 ;
        RECT 1.885 3.000 2.115 3.080 ;
        RECT 5.085 3.000 5.315 3.160 ;
        RECT 1.885 2.770 5.315 3.000 ;
        RECT 6.685 2.970 6.915 3.160 ;
        RECT 1.885 2.695 2.115 2.770 ;
        RECT 2.325 2.310 4.770 2.540 ;
        RECT 2.325 1.955 2.555 2.310 ;
        RECT 2.135 1.945 2.555 1.955 ;
        RECT 1.245 1.595 2.555 1.945 ;
        RECT 1.245 0.985 1.475 1.595 ;
        RECT 2.135 1.590 2.555 1.595 ;
        RECT 4.540 1.930 4.770 2.310 ;
        RECT 4.540 1.570 4.945 1.930 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi21b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi21b_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi21b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.760 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 11.760 4.220 ;
        RECT 4.205 3.230 4.435 3.620 ;
        RECT 5.805 3.230 6.035 3.620 ;
        RECT 7.405 3.230 7.635 3.620 ;
        RECT 9.005 3.230 9.235 3.620 ;
        RECT 11.265 2.235 11.495 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 12.190 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 12.190 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 8.205 0.300 8.435 0.690 ;
        RECT 9.805 0.300 10.035 1.370 ;
        RECT 11.265 0.300 11.495 1.370 ;
        RECT 0.000 -0.300 11.760 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.515200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.935 2.265 3.095 2.495 ;
        RECT 2.750 1.275 3.095 2.265 ;
        RECT 0.805 1.045 6.895 1.275 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.380 1.590 2.520 1.955 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 10.935 1.600 11.335 1.965 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.580 1.590 7.260 1.955 ;
    END
  END B
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.105 3.690 3.335 ;
        RECT 0.205 2.870 0.435 3.105 ;
        RECT 3.460 3.000 3.690 3.105 ;
        RECT 9.805 3.000 10.035 3.300 ;
        RECT 3.460 2.770 10.035 3.000 ;
        RECT 3.760 2.310 8.010 2.540 ;
        RECT 3.760 1.955 3.990 2.310 ;
        RECT 3.565 1.590 3.990 1.955 ;
        RECT 7.780 1.955 8.010 2.310 ;
        RECT 7.780 1.915 9.660 1.955 ;
        RECT 10.465 1.915 10.695 3.390 ;
        RECT 7.780 1.650 10.695 1.915 ;
        RECT 7.780 1.590 9.660 1.650 ;
        RECT 7.405 0.990 9.235 1.220 ;
        RECT 10.465 0.990 10.695 1.650 ;
        RECT 7.405 0.760 7.635 0.990 ;
        RECT 4.100 0.530 7.635 0.760 ;
        RECT 9.005 0.655 9.235 0.990 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi21b_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi22_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi22_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 4.880 3.230 5.110 3.620 ;
        RECT 6.480 3.230 6.710 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 6.480 0.300 6.710 0.690 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.972000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 2.650 0.435 2.815 ;
        RECT 1.775 2.650 3.720 2.880 ;
        RECT 0.205 2.420 2.065 2.650 ;
        RECT 3.405 2.480 3.720 2.650 ;
        RECT 3.490 2.335 3.720 2.480 ;
        RECT 3.490 1.240 3.930 2.335 ;
        RECT 2.470 1.010 5.190 1.240 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 1.590 1.640 1.965 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.180 1.590 3.260 1.965 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.455 1.590 5.535 1.965 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 6.055 1.590 7.135 1.965 ;
    END
  END D
  OBS
      LAYER Metal1 ;
        RECT 0.935 3.160 4.310 3.390 ;
        RECT 4.080 2.765 4.310 3.160 ;
        RECT 7.280 2.765 7.510 2.885 ;
        RECT 4.080 2.535 7.510 2.765 ;
        RECT 0.205 1.000 2.035 1.230 ;
        RECT 0.205 0.535 0.435 1.000 ;
        RECT 1.805 0.760 2.035 1.000 ;
        RECT 5.680 1.010 7.565 1.240 ;
        RECT 5.680 0.780 5.910 1.010 ;
        RECT 1.805 0.530 3.690 0.760 ;
        RECT 4.015 0.550 5.910 0.780 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi22_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi22_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi22_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 8.045 3.230 8.275 3.620 ;
        RECT 9.645 3.230 9.875 3.620 ;
        RECT 11.245 3.230 11.475 3.620 ;
        RECT 12.845 3.230 13.075 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 11.245 0.300 11.475 0.690 ;
        RECT 12.845 0.300 13.075 0.690 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.950400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.915 2.700 6.135 2.930 ;
        RECT 4.070 1.220 4.435 2.700 ;
        RECT 4.070 0.990 9.940 1.220 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.490 1.625 3.260 1.920 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.665 1.600 6.460 1.960 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 7.620 1.630 10.390 1.925 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.820 1.630 13.500 1.925 ;
    END
  END D
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.160 6.890 3.390 ;
        RECT 0.205 2.200 0.435 3.160 ;
        RECT 6.605 2.930 6.835 3.160 ;
        RECT 13.645 2.930 13.875 3.390 ;
        RECT 6.605 2.700 13.875 2.930 ;
        RECT 6.605 2.635 6.835 2.700 ;
        RECT 13.645 2.235 13.875 2.700 ;
        RECT 0.205 1.150 0.435 1.185 ;
        RECT 0.205 0.920 3.635 1.150 ;
        RECT 0.205 0.740 0.435 0.920 ;
        RECT 3.405 0.760 3.635 0.920 ;
        RECT 10.445 0.990 13.875 1.220 ;
        RECT 10.445 0.760 10.675 0.990 ;
        RECT 13.645 0.795 13.875 0.990 ;
        RECT 3.405 0.530 6.895 0.760 ;
        RECT 7.160 0.530 10.675 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi22_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi31_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi31_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.845 3.230 5.075 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 6.450 0.300 6.680 0.690 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 1.630 1.660 1.925 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.180 1.630 3.260 1.925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.420 1.630 5.500 1.925 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.124500 ;
    PORT
      LAYER Metal1 ;
        RECT 6.355 2.320 7.015 2.550 ;
        RECT 6.730 1.220 7.015 2.320 ;
        RECT 5.645 0.990 7.535 1.220 ;
        RECT 5.645 0.760 5.875 0.990 ;
        RECT 3.970 0.530 5.875 0.760 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 5.910 1.630 6.500 1.925 ;
    END
  END D
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.950 0.435 3.390 ;
        RECT 1.805 2.950 2.035 3.390 ;
        RECT 3.405 2.950 3.635 3.390 ;
        RECT 3.910 2.950 4.140 3.390 ;
        RECT 5.645 3.160 7.480 3.390 ;
        RECT 5.645 2.950 5.875 3.160 ;
        RECT 0.205 2.720 5.875 2.950 ;
        RECT 0.205 2.200 0.435 2.720 ;
        RECT 1.805 2.200 2.035 2.720 ;
        RECT 3.405 2.200 3.635 2.720 ;
        RECT 3.910 2.200 4.140 2.720 ;
        RECT 5.645 2.200 5.875 2.720 ;
        RECT 7.250 2.200 7.480 3.160 ;
        RECT 0.205 1.150 0.435 1.170 ;
        RECT 0.205 0.920 2.035 1.150 ;
        RECT 2.470 0.990 5.130 1.220 ;
        RECT 0.205 0.800 0.435 0.920 ;
        RECT 1.805 0.760 2.035 0.920 ;
        RECT 1.805 0.530 3.695 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi31_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__aoi31_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__aoi31_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.560 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.205 3.230 4.435 3.620 ;
        RECT 5.805 3.230 6.035 3.620 ;
        RECT 8.045 3.230 8.275 3.620 ;
        RECT 9.645 3.230 9.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.990 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 11.245 0.300 11.475 0.690 ;
        RECT 12.845 0.300 13.075 0.690 ;
        RECT 0.000 -0.300 14.560 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.470 1.615 3.265 1.925 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.780 1.590 6.460 1.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 7.620 1.590 10.300 1.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 10.820 1.590 13.495 1.950 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.875200 ;
    PORT
      LAYER Metal1 ;
        RECT 11.185 2.700 14.070 2.930 ;
        RECT 13.725 1.220 14.070 2.700 ;
        RECT 7.155 0.990 14.070 1.220 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.940 0.435 3.390 ;
        RECT 1.805 2.940 2.035 3.390 ;
        RECT 3.405 2.940 3.635 3.390 ;
        RECT 5.005 2.940 5.235 3.390 ;
        RECT 6.605 2.940 6.835 3.390 ;
        RECT 8.845 2.940 9.075 3.390 ;
        RECT 10.350 3.160 13.930 3.390 ;
        RECT 10.350 2.940 10.580 3.160 ;
        RECT 0.205 2.710 10.580 2.940 ;
        RECT 0.205 2.200 0.435 2.710 ;
        RECT 1.805 2.200 2.035 2.710 ;
        RECT 3.405 2.200 3.635 2.710 ;
        RECT 5.005 2.200 5.235 2.710 ;
        RECT 6.605 2.200 6.835 2.710 ;
        RECT 8.845 2.200 9.075 2.710 ;
        RECT 3.400 1.150 6.890 1.220 ;
        RECT 0.205 0.990 6.890 1.150 ;
        RECT 0.205 0.920 3.700 0.990 ;
        RECT 0.205 0.530 0.435 0.920 ;
        RECT 4.070 0.530 9.930 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__aoi31_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_12
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 0.205 2.850 0.435 3.620 ;
        RECT 1.805 2.765 2.035 3.620 ;
        RECT 3.405 2.770 3.635 3.620 ;
        RECT 5.005 2.770 5.235 3.620 ;
        RECT 6.605 2.765 6.835 3.620 ;
        RECT 8.205 2.265 8.435 3.620 ;
        RECT 9.820 2.265 10.050 3.620 ;
        RECT 11.420 2.265 11.650 3.620 ;
        RECT 13.020 2.265 13.250 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.840 ;
        RECT 1.805 0.300 2.035 0.710 ;
        RECT 3.405 0.300 3.635 0.710 ;
        RECT 5.005 0.300 5.235 0.710 ;
        RECT 6.605 0.300 6.835 0.710 ;
        RECT 8.205 0.300 8.435 1.300 ;
        RECT 9.820 0.300 10.050 1.300 ;
        RECT 11.420 0.300 11.650 1.300 ;
        RECT 13.020 0.300 13.250 1.300 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 1.570 3.145 2.075 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.461300 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 2.535 4.435 3.390 ;
        RECT 5.805 2.535 6.035 3.390 ;
        RECT 7.405 2.535 7.635 3.390 ;
        RECT 4.205 2.305 7.635 2.535 ;
        RECT 7.405 2.035 7.635 2.305 ;
        RECT 9.020 2.035 9.250 3.390 ;
        RECT 10.620 2.035 10.850 3.390 ;
        RECT 12.220 2.035 12.450 3.390 ;
        RECT 7.405 1.530 12.450 2.035 ;
        RECT 7.405 1.330 7.635 1.530 ;
        RECT 4.205 1.100 7.635 1.330 ;
        RECT 4.205 0.990 4.435 1.100 ;
        RECT 5.805 0.990 6.035 1.100 ;
        RECT 7.405 0.990 7.635 1.100 ;
        RECT 9.020 0.990 9.250 1.530 ;
        RECT 10.620 0.990 10.850 1.530 ;
        RECT 12.220 0.990 12.450 1.530 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.535 1.235 3.390 ;
        RECT 2.605 2.535 2.835 3.390 ;
        RECT 1.005 2.305 3.605 2.535 ;
        RECT 3.375 1.920 3.605 2.305 ;
        RECT 3.375 1.630 7.175 1.920 ;
        RECT 3.375 1.330 3.605 1.630 ;
        RECT 1.005 1.100 3.605 1.330 ;
        RECT 1.005 0.990 1.235 1.100 ;
        RECT 2.605 0.990 2.835 1.100 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_12


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.660 2.265 2.890 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 3.790 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 3.790 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.660 0.300 2.890 1.400 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.570 0.675 2.285 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 0.530 2.200 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.895 0.435 3.380 ;
        RECT 0.205 2.665 1.330 2.895 ;
        RECT 1.100 2.030 1.330 2.665 ;
        RECT 1.100 1.575 1.395 2.030 ;
        RECT 1.100 1.175 1.330 1.575 ;
        RECT 0.205 0.945 1.330 1.175 ;
        RECT 0.205 0.795 0.435 0.945 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.205 2.140 4.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 4.205 0.300 4.435 1.370 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.570 0.675 2.285 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 2.040 2.200 3.390 ;
        RECT 3.405 2.040 3.800 3.390 ;
        RECT 1.805 1.755 3.800 2.040 ;
        RECT 1.805 0.530 2.200 1.755 ;
        RECT 3.405 0.530 3.800 1.755 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.895 0.435 3.380 ;
        RECT 0.205 2.665 1.330 2.895 ;
        RECT 1.100 2.030 1.330 2.665 ;
        RECT 1.100 1.575 1.395 2.030 ;
        RECT 1.100 1.175 1.330 1.575 ;
        RECT 0.205 0.945 1.330 1.175 ;
        RECT 0.205 0.795 0.435 0.945 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__buff_8
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__buff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.205 3.185 0.435 3.620 ;
        RECT 1.805 2.265 2.035 3.620 ;
        RECT 3.405 2.180 3.635 3.620 ;
        RECT 5.005 2.210 5.235 3.620 ;
        RECT 6.605 2.210 6.835 3.620 ;
        RECT 8.205 2.210 8.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.735 ;
        RECT 1.805 0.300 2.035 1.275 ;
        RECT 3.405 0.300 3.635 1.370 ;
        RECT 5.005 0.300 5.235 1.340 ;
        RECT 6.605 0.300 6.835 1.340 ;
        RECT 8.205 0.300 8.435 1.325 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 2.060 0.585 2.405 ;
        RECT 0.205 1.610 0.770 2.060 ;
        RECT 0.205 1.455 0.585 1.610 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.283200 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 1.980 4.435 3.390 ;
        RECT 5.805 1.980 6.035 3.390 ;
        RECT 7.405 1.980 7.635 3.390 ;
        RECT 9.005 1.980 9.235 3.390 ;
        RECT 4.205 1.570 9.235 1.980 ;
        RECT 4.205 0.990 4.435 1.570 ;
        RECT 5.805 0.990 6.035 1.570 ;
        RECT 7.405 0.990 7.635 1.570 ;
        RECT 9.005 0.990 9.235 1.570 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.035 1.235 3.390 ;
        RECT 2.605 2.035 2.835 3.390 ;
        RECT 1.005 1.995 2.835 2.035 ;
        RECT 1.005 1.935 3.065 1.995 ;
        RECT 1.005 1.805 3.975 1.935 ;
        RECT 1.005 0.990 1.235 1.805 ;
        RECT 2.605 1.660 3.975 1.805 ;
        RECT 2.605 1.610 3.065 1.660 ;
        RECT 2.605 0.990 2.835 1.610 ;
  END
END gf180mcu_as_sc_mcu7t3v3__buff_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__clkbuff_12
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__clkbuff_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 14.000 4.220 ;
        RECT 0.205 2.850 0.435 3.620 ;
        RECT 1.805 2.765 2.035 3.620 ;
        RECT 3.405 2.770 3.635 3.620 ;
        RECT 5.005 2.770 5.235 3.620 ;
        RECT 6.605 2.765 6.835 3.620 ;
        RECT 8.205 2.265 8.435 3.620 ;
        RECT 9.820 2.265 10.050 3.620 ;
        RECT 11.420 2.265 11.650 3.620 ;
        RECT 13.020 2.265 13.250 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 14.430 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 14.430 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.700 ;
        RECT 1.805 0.300 2.035 0.710 ;
        RECT 3.405 0.300 3.635 0.710 ;
        RECT 5.005 0.300 5.235 0.710 ;
        RECT 6.605 0.300 6.835 0.710 ;
        RECT 8.205 0.300 8.435 0.690 ;
        RECT 9.820 0.300 10.050 0.690 ;
        RECT 11.420 0.300 11.650 0.690 ;
        RECT 13.020 0.300 13.250 0.690 ;
        RECT 0.000 -0.300 14.000 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.515 1.570 3.145 2.075 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 2.535 4.435 3.390 ;
        RECT 5.805 2.535 6.035 3.390 ;
        RECT 7.405 2.535 7.635 3.390 ;
        RECT 4.205 2.305 7.635 2.535 ;
        RECT 7.405 2.035 7.635 2.305 ;
        RECT 9.020 2.035 9.250 3.390 ;
        RECT 10.620 2.035 10.850 3.390 ;
        RECT 12.220 2.035 12.450 3.390 ;
        RECT 7.405 1.530 12.450 2.035 ;
        RECT 7.405 1.330 7.635 1.530 ;
        RECT 4.205 1.100 7.635 1.330 ;
        RECT 4.205 0.530 4.435 1.100 ;
        RECT 5.805 0.530 6.035 1.100 ;
        RECT 7.405 0.530 7.635 1.100 ;
        RECT 9.020 0.530 9.250 1.530 ;
        RECT 10.620 0.530 10.850 1.530 ;
        RECT 12.220 0.530 12.450 1.530 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.535 1.235 3.390 ;
        RECT 2.605 2.535 2.835 3.390 ;
        RECT 1.005 2.305 3.605 2.535 ;
        RECT 3.375 1.920 3.605 2.305 ;
        RECT 3.375 1.630 7.175 1.920 ;
        RECT 3.375 1.330 3.605 1.630 ;
        RECT 1.005 1.100 3.605 1.330 ;
        RECT 1.005 0.530 1.235 1.100 ;
        RECT 2.605 0.530 2.835 1.100 ;
  END
END gf180mcu_as_sc_mcu7t3v3__clkbuff_12


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__clkbuff_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__clkbuff_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.040 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.040 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
        RECT 4.205 2.140 4.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 5.470 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 5.470 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 4.205 0.300 4.435 0.730 ;
        RECT 0.000 -0.300 5.040 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.570 0.675 2.285 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.184000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.805 2.040 2.200 3.390 ;
        RECT 3.405 2.040 3.800 3.390 ;
        RECT 1.805 1.755 3.800 2.040 ;
        RECT 1.805 0.530 2.200 1.755 ;
        RECT 3.405 0.530 3.800 1.755 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.895 0.435 3.380 ;
        RECT 0.205 2.665 1.330 2.895 ;
        RECT 1.100 2.030 1.330 2.665 ;
        RECT 1.100 1.575 1.395 2.030 ;
        RECT 1.100 1.175 1.330 1.575 ;
        RECT 0.205 0.945 1.330 1.175 ;
        RECT 0.205 0.530 0.435 0.945 ;
  END
END gf180mcu_as_sc_mcu7t3v3__clkbuff_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__clkbuff_8
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__clkbuff_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 10.080 4.220 ;
        RECT 0.205 3.185 0.435 3.620 ;
        RECT 1.805 2.265 2.035 3.620 ;
        RECT 3.405 2.180 3.635 3.620 ;
        RECT 5.005 2.210 5.235 3.620 ;
        RECT 6.605 2.210 6.835 3.620 ;
        RECT 8.205 2.210 8.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 10.510 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 10.510 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.735 ;
        RECT 1.805 0.300 2.035 0.700 ;
        RECT 3.405 0.300 3.635 0.795 ;
        RECT 5.005 0.300 5.235 0.765 ;
        RECT 6.605 0.300 6.835 0.765 ;
        RECT 8.205 0.300 8.435 0.750 ;
        RECT 0.000 -0.300 10.080 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.764000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 2.060 0.585 2.405 ;
        RECT 0.205 1.610 0.770 2.060 ;
        RECT 0.205 1.455 0.585 1.610 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.544000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.205 1.980 4.435 3.390 ;
        RECT 5.805 1.980 6.035 3.390 ;
        RECT 7.405 1.980 7.635 3.390 ;
        RECT 9.005 1.980 9.235 3.390 ;
        RECT 4.205 1.570 9.235 1.980 ;
        RECT 4.205 0.710 4.435 1.570 ;
        RECT 5.805 0.710 6.035 1.570 ;
        RECT 7.405 0.710 7.635 1.570 ;
        RECT 9.005 0.710 9.235 1.570 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.005 2.035 1.235 3.390 ;
        RECT 2.605 2.035 2.835 3.390 ;
        RECT 1.005 1.995 2.835 2.035 ;
        RECT 1.005 1.935 3.065 1.995 ;
        RECT 1.005 1.805 3.975 1.935 ;
        RECT 1.005 0.710 1.235 1.805 ;
        RECT 2.605 1.660 3.975 1.805 ;
        RECT 2.605 1.610 3.065 1.660 ;
        RECT 2.605 0.710 2.835 1.610 ;
  END
END gf180mcu_as_sc_mcu7t3v3__clkbuff_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__dfsrtp_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__dfsrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 20.720 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.490 3.230 2.720 3.620 ;
        RECT 7.120 3.285 7.540 3.620 ;
        RECT 9.480 3.285 9.845 3.620 ;
        RECT 14.085 3.200 14.315 3.620 ;
        RECT 15.930 3.210 16.160 3.620 ;
        RECT 17.860 2.145 18.090 3.620 ;
        RECT 18.510 2.145 18.740 3.620 ;
        RECT 20.110 2.145 20.340 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 21.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 21.150 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.490 0.300 2.720 0.690 ;
        RECT 8.195 0.300 8.550 0.635 ;
        RECT 15.900 0.300 16.315 0.635 ;
        RECT 18.510 0.300 18.740 1.390 ;
        RECT 20.110 0.300 20.340 1.385 ;
        RECT 0.000 -0.300 20.720 0.300 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 1.600 0.860 2.060 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 19.215 0.530 19.645 3.390 ;
    END
  END Q
  PIN RN
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 7.595 1.560 8.730 1.790 ;
        RECT 8.500 1.295 8.730 1.560 ;
        RECT 8.500 1.065 9.735 1.295 ;
        RECT 15.955 1.115 16.620 1.990 ;
        RECT 9.505 0.760 9.735 1.065 ;
        RECT 15.435 0.880 16.620 1.115 ;
        RECT 15.435 0.760 15.670 0.880 ;
        RECT 9.505 0.530 15.670 0.760 ;
    END
  END RN
  PIN SN
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 10.075 2.835 11.910 3.040 ;
        RECT 10.075 2.810 11.925 2.835 ;
        RECT 10.075 1.625 10.305 2.810 ;
        RECT 11.650 2.570 11.925 2.810 ;
        RECT 11.650 2.520 11.910 2.570 ;
        RECT 13.575 1.565 14.725 2.510 ;
      LAYER Metal2 ;
        RECT 11.635 2.560 11.925 2.900 ;
        RECT 11.645 1.960 11.925 2.560 ;
        RECT 11.645 1.680 13.965 1.960 ;
    END
  END SN
  PIN D
    ANTENNAGATEAREA 0.673300 ;
    PORT
      LAYER Metal1 ;
        RECT 2.345 1.400 3.180 2.535 ;
    END
  END D
  OBS
      LAYER Metal1 ;
        RECT 3.000 3.160 5.620 3.390 ;
        RECT 3.000 3.000 3.230 3.160 ;
        RECT 0.205 2.935 0.445 2.995 ;
        RECT 1.105 2.935 3.230 3.000 ;
        RECT 0.205 2.770 3.230 2.935 ;
        RECT 0.205 2.705 1.335 2.770 ;
        RECT 0.205 2.650 0.445 2.705 ;
        RECT 1.105 1.985 1.335 2.705 ;
        RECT 3.465 2.530 3.695 2.925 ;
        RECT 4.470 2.575 4.700 3.160 ;
        RECT 1.745 2.265 2.095 2.495 ;
        RECT 3.410 2.285 3.695 2.530 ;
        RECT 1.105 1.605 1.405 1.985 ;
        RECT 0.205 1.275 0.435 1.330 ;
        RECT 1.105 1.275 1.335 1.605 ;
        RECT 0.205 1.045 1.335 1.275 ;
        RECT 1.805 1.170 2.035 2.265 ;
        RECT 0.205 0.990 0.435 1.045 ;
        RECT 1.800 0.940 3.180 1.170 ;
        RECT 3.410 0.990 3.640 2.285 ;
        RECT 4.440 2.195 4.700 2.575 ;
        RECT 2.950 0.760 3.180 0.940 ;
        RECT 3.870 0.760 4.100 2.100 ;
        RECT 4.470 1.570 4.700 2.195 ;
        RECT 4.930 1.365 5.160 2.900 ;
        RECT 5.390 1.630 5.620 3.160 ;
        RECT 5.910 3.055 6.140 3.170 ;
        RECT 8.005 3.055 8.235 3.180 ;
        RECT 5.910 2.825 8.235 3.055 ;
        RECT 8.660 3.055 8.890 3.165 ;
        RECT 8.660 2.825 9.830 3.055 ;
        RECT 5.850 2.365 9.285 2.595 ;
        RECT 5.850 1.365 6.080 2.365 ;
        RECT 9.055 2.025 9.285 2.365 ;
        RECT 4.930 1.135 6.080 1.365 ;
        RECT 6.315 1.315 6.545 1.835 ;
        RECT 6.835 1.560 7.220 2.015 ;
        RECT 9.035 1.560 9.355 2.025 ;
        RECT 9.600 2.015 9.830 2.825 ;
        RECT 12.155 2.970 12.385 3.390 ;
        RECT 14.545 3.150 15.700 3.380 ;
        RECT 14.545 2.970 14.775 3.150 ;
        RECT 12.155 2.740 14.775 2.970 ;
        RECT 15.470 2.965 15.700 3.150 ;
        RECT 16.390 3.160 17.540 3.390 ;
        RECT 16.390 2.965 16.620 3.160 ;
        RECT 9.585 1.635 9.845 2.015 ;
        RECT 7.170 1.315 7.550 1.330 ;
        RECT 4.930 0.990 5.160 1.135 ;
        RECT 6.315 1.085 7.550 1.315 ;
        RECT 10.535 1.275 10.795 2.550 ;
        RECT 11.025 2.290 11.285 2.580 ;
        RECT 11.025 2.030 11.925 2.290 ;
        RECT 6.315 0.760 6.545 1.085 ;
        RECT 7.170 1.070 7.550 1.085 ;
        RECT 10.435 1.045 10.795 1.275 ;
        RECT 11.030 0.990 11.290 1.800 ;
        RECT 11.695 1.625 11.925 2.030 ;
        RECT 12.155 1.275 12.385 2.740 ;
        RECT 13.000 2.275 13.340 2.505 ;
        RECT 11.520 1.045 12.385 1.275 ;
        RECT 12.620 1.390 12.850 2.080 ;
        RECT 12.620 1.010 12.880 1.390 ;
        RECT 13.110 1.325 13.340 2.275 ;
        RECT 15.005 1.920 15.235 2.920 ;
        RECT 15.470 2.735 16.620 2.965 ;
        RECT 16.850 2.465 17.080 2.925 ;
        RECT 14.970 1.665 15.235 1.920 ;
        RECT 15.465 2.235 17.080 2.465 ;
        RECT 14.970 1.325 15.200 1.665 ;
        RECT 15.465 1.615 15.695 2.235 ;
        RECT 16.850 1.575 17.080 2.235 ;
        RECT 17.310 2.035 17.540 3.160 ;
        RECT 17.310 1.805 17.650 2.035 ;
        RECT 18.050 1.685 18.955 1.915 ;
        RECT 18.050 1.575 18.280 1.685 ;
        RECT 16.850 1.345 18.280 1.575 ;
        RECT 13.110 1.045 15.200 1.325 ;
        RECT 2.950 0.530 6.545 0.760 ;
        RECT 17.770 0.705 18.000 1.345 ;
      LAYER Metal2 ;
        RECT 4.380 2.245 11.350 2.530 ;
        RECT 6.830 1.680 10.855 1.965 ;
        RECT 7.170 1.060 12.945 1.340 ;
        RECT 7.170 1.055 7.510 1.060 ;
  END
END gf180mcu_as_sc_mcu7t3v3__dfsrtp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__dfxtn_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__dfxtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.490 3.230 2.720 3.620 ;
        RECT 7.000 3.230 7.230 3.620 ;
        RECT 11.360 3.230 11.590 3.620 ;
        RECT 12.910 2.145 13.140 3.620 ;
        RECT 14.510 2.145 14.740 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 15.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.490 0.300 2.720 0.690 ;
        RECT 7.000 0.300 7.230 0.690 ;
        RECT 11.360 0.300 11.590 0.690 ;
        RECT 12.910 0.300 13.140 1.390 ;
        RECT 14.510 0.300 14.740 1.385 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 1.600 0.860 2.060 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.985 1.630 4.430 2.930 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.615 0.990 14.045 2.550 ;
    END
  END Q
  OBS
      LAYER Metal1 ;
        RECT 1.790 3.000 2.035 3.390 ;
        RECT 2.970 3.160 6.205 3.390 ;
        RECT 2.970 3.000 3.200 3.160 ;
        RECT 0.205 2.935 0.445 2.995 ;
        RECT 0.205 2.705 1.335 2.935 ;
        RECT 0.205 2.650 0.445 2.705 ;
        RECT 1.105 1.985 1.335 2.705 ;
        RECT 1.790 2.770 3.200 3.000 ;
        RECT 1.790 2.450 2.035 2.770 ;
        RECT 1.105 1.605 1.405 1.985 ;
        RECT 0.205 1.275 0.435 1.330 ;
        RECT 1.105 1.275 1.335 1.605 ;
        RECT 1.790 1.550 2.020 2.450 ;
        RECT 2.250 2.045 3.680 2.275 ;
        RECT 2.250 1.720 2.480 2.045 ;
        RECT 1.790 1.280 2.035 1.550 ;
        RECT 2.850 1.280 3.080 1.790 ;
        RECT 0.205 1.045 1.335 1.275 ;
        RECT 1.750 1.045 3.080 1.280 ;
        RECT 0.205 0.990 0.435 1.045 ;
        RECT 3.450 0.760 3.680 2.045 ;
        RECT 4.660 1.400 4.890 2.550 ;
        RECT 5.120 1.630 5.350 3.160 ;
        RECT 5.925 3.090 6.205 3.160 ;
        RECT 5.925 2.755 6.305 3.090 ;
        RECT 8.320 3.005 10.620 3.235 ;
        RECT 5.580 2.295 7.530 2.525 ;
        RECT 5.580 1.400 5.810 2.295 ;
        RECT 6.045 1.990 6.325 2.025 ;
        RECT 4.660 1.170 5.810 1.400 ;
        RECT 6.040 1.645 6.325 1.990 ;
        RECT 4.660 0.990 4.890 1.170 ;
        RECT 6.040 0.760 6.270 1.645 ;
        RECT 6.625 1.640 6.885 1.990 ;
        RECT 6.655 1.220 6.885 1.640 ;
        RECT 7.300 1.625 7.530 2.295 ;
        RECT 7.800 1.220 8.030 2.550 ;
        RECT 8.320 1.985 8.550 3.005 ;
        RECT 8.260 1.595 8.640 1.985 ;
        RECT 8.870 1.560 9.190 2.025 ;
        RECT 6.655 0.990 8.030 1.220 ;
        RECT 9.420 1.150 9.650 2.550 ;
        RECT 10.390 1.625 10.620 3.005 ;
        RECT 12.270 2.500 12.500 3.390 ;
        RECT 11.010 2.270 12.500 2.500 ;
        RECT 11.010 1.625 11.240 2.270 ;
        RECT 12.270 1.980 12.500 2.270 ;
        RECT 11.810 1.150 12.040 1.980 ;
        RECT 9.420 0.920 12.040 1.150 ;
        RECT 12.270 1.620 12.650 1.980 ;
        RECT 12.270 0.990 12.500 1.620 ;
        RECT 3.450 0.530 6.270 0.760 ;
      LAYER Metal2 ;
        RECT 5.915 2.760 9.200 3.040 ;
        RECT 6.045 1.975 6.325 2.025 ;
        RECT 6.035 1.695 8.640 1.975 ;
        RECT 6.045 1.645 6.325 1.695 ;
        RECT 8.920 1.640 9.200 2.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__dfxtn_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__dfxtp_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 15.120 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.490 3.230 2.720 3.620 ;
        RECT 7.000 3.230 7.230 3.620 ;
        RECT 11.360 3.230 11.590 3.620 ;
        RECT 12.910 2.145 13.140 3.620 ;
        RECT 14.510 2.145 14.740 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 15.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 15.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.490 0.300 2.720 0.690 ;
        RECT 7.000 0.300 7.230 0.690 ;
        RECT 11.360 0.300 11.590 0.690 ;
        RECT 12.910 0.300 13.140 1.390 ;
        RECT 14.510 0.300 14.740 1.385 ;
        RECT 0.000 -0.300 15.120 0.300 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.125 1.600 0.860 2.060 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.985 1.630 4.430 2.930 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 13.615 0.990 14.045 2.550 ;
    END
  END Q
  OBS
      LAYER Metal1 ;
        RECT 2.970 3.160 6.205 3.390 ;
        RECT 2.970 3.000 3.200 3.160 ;
        RECT 0.205 2.935 0.445 2.995 ;
        RECT 1.105 2.935 3.200 3.000 ;
        RECT 0.205 2.770 3.200 2.935 ;
        RECT 0.205 2.705 1.335 2.770 ;
        RECT 0.205 2.650 0.445 2.705 ;
        RECT 1.105 1.985 1.335 2.705 ;
        RECT 1.745 2.265 2.095 2.495 ;
        RECT 1.805 2.000 2.035 2.265 ;
        RECT 1.105 1.605 1.405 1.985 ;
        RECT 1.805 1.770 3.680 2.000 ;
        RECT 0.205 1.275 0.435 1.330 ;
        RECT 1.105 1.275 1.335 1.605 ;
        RECT 0.205 1.045 1.335 1.275 ;
        RECT 0.205 0.990 0.435 1.045 ;
        RECT 1.805 0.990 2.035 1.770 ;
        RECT 3.375 1.640 3.680 1.770 ;
        RECT 3.450 0.760 3.680 1.640 ;
        RECT 4.660 1.400 4.890 2.550 ;
        RECT 5.120 1.630 5.350 3.160 ;
        RECT 5.925 3.090 6.205 3.160 ;
        RECT 5.925 2.755 6.305 3.090 ;
        RECT 8.320 3.005 10.620 3.235 ;
        RECT 5.580 2.295 7.530 2.525 ;
        RECT 5.580 1.400 5.810 2.295 ;
        RECT 6.045 1.990 6.325 2.025 ;
        RECT 4.660 1.170 5.810 1.400 ;
        RECT 6.040 1.645 6.325 1.990 ;
        RECT 4.660 0.990 4.890 1.170 ;
        RECT 6.040 0.760 6.270 1.645 ;
        RECT 6.625 1.640 6.885 1.990 ;
        RECT 6.655 1.220 6.885 1.640 ;
        RECT 7.300 1.625 7.530 2.295 ;
        RECT 7.800 1.220 8.030 2.550 ;
        RECT 8.320 1.985 8.550 3.005 ;
        RECT 8.260 1.595 8.640 1.985 ;
        RECT 8.870 1.560 9.190 2.025 ;
        RECT 6.655 0.990 8.030 1.220 ;
        RECT 9.420 1.150 9.650 2.550 ;
        RECT 10.390 1.625 10.620 3.005 ;
        RECT 12.270 2.500 12.500 3.390 ;
        RECT 11.010 2.270 12.500 2.500 ;
        RECT 11.010 1.625 11.240 2.270 ;
        RECT 12.270 1.980 12.500 2.270 ;
        RECT 11.810 1.150 12.040 1.980 ;
        RECT 9.420 0.920 12.040 1.150 ;
        RECT 12.270 1.620 12.650 1.980 ;
        RECT 12.270 0.990 12.500 1.620 ;
        RECT 3.450 0.530 6.270 0.760 ;
      LAYER Metal2 ;
        RECT 5.915 2.760 9.200 3.040 ;
        RECT 6.045 1.975 6.325 2.025 ;
        RECT 6.035 1.695 8.640 1.975 ;
        RECT 6.045 1.645 6.325 1.695 ;
        RECT 8.920 1.640 9.200 2.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__dfxtp_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 1.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal1 ;
        RECT 0.330 0.805 0.630 2.750 ;
    END
  END DIODE
END gf180mcu_as_sc_mcu7t3v3__diode_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_1
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.560 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 0.560 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 0.990 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 0.990 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 0.560 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_1


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_2
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 1.550 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_4
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fill_8
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__fill_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fillcap_16
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fillcap_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 8.525 2.555 8.755 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.740 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.240 1.735 0.470 3.390 ;
        RECT 8.020 2.095 8.755 2.325 ;
        RECT 0.240 1.500 1.040 1.735 ;
        RECT 0.650 1.440 1.040 1.500 ;
        RECT 8.525 0.980 8.755 2.095 ;
  END
END gf180mcu_as_sc_mcu7t3v3__fillcap_16


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fillcap_4
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fillcap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 1.805 2.565 2.035 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.740 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.240 1.735 0.470 3.390 ;
        RECT 1.305 2.090 2.035 2.335 ;
        RECT 0.240 1.500 1.040 1.735 ;
        RECT 0.650 1.440 1.040 1.500 ;
        RECT 1.805 0.530 2.035 2.090 ;
  END
END gf180mcu_as_sc_mcu7t3v3__fillcap_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__fillcap_8
  CLASS CORE SPACER ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__fillcap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.480 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 4.480 4.220 ;
        RECT 4.045 2.565 4.275 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.910 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.910 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.740 ;
        RECT 0.000 -0.300 4.480 0.300 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 0.240 1.735 0.470 3.390 ;
        RECT 3.520 2.095 4.275 2.335 ;
        RECT 0.240 1.500 1.040 1.735 ;
        RECT 0.650 1.440 1.040 1.500 ;
        RECT 4.045 0.980 4.275 2.095 ;
  END
END gf180mcu_as_sc_mcu7t3v3__fillcap_8


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__inv_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.205 2.355 0.435 3.620 ;
        RECT 1.805 2.295 2.035 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.235 ;
        RECT 1.805 0.300 2.035 1.235 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.255 1.235 3.385 ;
        RECT 1.005 1.260 1.350 2.255 ;
        RECT 1.005 0.530 1.235 1.260 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.590 0.775 2.125 ;
    END
  END A
END gf180mcu_as_sc_mcu7t3v3__inv_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__inv_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 0.205 2.355 0.435 3.620 ;
        RECT 1.805 2.295 2.035 3.620 ;
        RECT 3.405 2.175 3.635 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.235 ;
        RECT 1.805 0.300 2.035 1.235 ;
        RECT 3.405 0.300 3.635 1.395 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.255 1.235 3.385 ;
        RECT 1.005 1.935 1.350 2.255 ;
        RECT 2.605 1.935 2.835 3.385 ;
        RECT 1.005 1.705 2.835 1.935 ;
        RECT 1.005 1.260 1.350 1.705 ;
        RECT 1.005 0.990 1.235 1.260 ;
        RECT 2.605 0.990 2.835 1.705 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.590 0.775 2.125 ;
    END
  END A
END gf180mcu_as_sc_mcu7t3v3__inv_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__inv_6
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__inv_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.205 2.355 0.435 3.620 ;
        RECT 1.805 2.295 2.035 3.620 ;
        RECT 3.405 2.175 3.635 3.620 ;
        RECT 5.005 2.175 5.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.235 ;
        RECT 1.805 0.300 2.035 1.235 ;
        RECT 3.405 0.300 3.635 1.395 ;
        RECT 5.005 0.300 5.235 1.395 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.712800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.255 1.235 3.385 ;
        RECT 1.005 1.935 1.350 2.255 ;
        RECT 2.605 1.935 2.835 3.385 ;
        RECT 4.205 1.935 4.570 3.385 ;
        RECT 1.005 1.705 4.570 1.935 ;
        RECT 1.005 1.260 1.350 1.705 ;
        RECT 1.005 0.990 1.235 1.260 ;
        RECT 2.605 0.990 2.835 1.705 ;
        RECT 4.205 0.990 4.570 1.705 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.998400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.590 0.775 2.125 ;
    END
  END A
END gf180mcu_as_sc_mcu7t3v3__inv_6


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__invz_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__invz_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 1.105 3.145 1.335 3.620 ;
        RECT 5.145 3.160 5.375 3.620 ;
        RECT 7.595 3.160 7.825 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.750 ;
        RECT 5.090 0.300 5.430 0.635 ;
        RECT 7.645 0.300 7.875 1.250 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  PIN EN
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.670 1.975 2.195 2.450 ;
        RECT 0.670 1.570 0.900 1.975 ;
        RECT 1.965 1.600 2.195 1.975 ;
    END
  END EN
  PIN A
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 7.135 2.050 8.190 2.450 ;
        RECT 7.960 1.650 8.190 2.050 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA 2.144600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.205 2.230 6.905 2.910 ;
        RECT 6.565 1.430 6.905 2.230 ;
        RECT 6.305 0.990 6.905 1.430 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.915 0.435 3.390 ;
        RECT 2.230 3.145 4.020 3.390 ;
        RECT 0.205 2.685 2.880 2.915 ;
        RECT 0.205 1.335 0.435 2.685 ;
        RECT 2.650 2.090 2.880 2.685 ;
        RECT 3.125 2.510 3.355 2.900 ;
        RECT 3.125 2.265 3.425 2.510 ;
        RECT 2.650 1.750 2.965 2.090 ;
        RECT 1.290 1.515 1.630 1.745 ;
        RECT 3.195 1.590 3.425 2.265 ;
        RECT 1.290 1.335 1.575 1.515 ;
        RECT 0.205 1.100 1.575 1.335 ;
        RECT 3.155 1.360 3.425 1.590 ;
        RECT 3.790 1.565 4.020 3.145 ;
        RECT 5.685 3.150 7.365 3.380 ;
        RECT 5.685 2.840 5.915 3.150 ;
        RECT 4.360 2.610 5.915 2.840 ;
        RECT 7.135 2.915 7.365 3.150 ;
        RECT 8.445 2.915 8.675 3.390 ;
        RECT 7.135 2.685 8.675 2.915 ;
        RECT 4.360 2.035 4.590 2.610 ;
        RECT 4.250 1.805 4.590 2.035 ;
        RECT 4.825 2.150 5.975 2.380 ;
        RECT 4.825 1.565 5.055 2.150 ;
        RECT 5.745 2.000 5.975 2.150 ;
        RECT 0.205 0.945 0.435 1.100 ;
        RECT 1.805 0.760 2.035 1.290 ;
        RECT 3.155 0.760 3.385 1.360 ;
        RECT 3.790 1.335 5.055 1.565 ;
        RECT 3.790 1.235 4.020 1.335 ;
        RECT 3.620 0.990 4.020 1.235 ;
        RECT 5.285 1.105 5.515 1.845 ;
        RECT 5.745 1.710 6.335 2.000 ;
        RECT 6.105 1.660 6.335 1.710 ;
        RECT 7.185 1.480 7.575 1.820 ;
        RECT 4.615 0.865 6.060 1.105 ;
        RECT 4.615 0.760 4.855 0.865 ;
        RECT 1.805 0.530 4.855 0.760 ;
        RECT 5.830 0.760 6.060 0.865 ;
        RECT 7.185 0.760 7.415 1.480 ;
        RECT 8.445 0.945 8.675 2.685 ;
        RECT 5.830 0.530 7.415 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__invz_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__maj3_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__maj3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 1.525 3.230 1.755 3.620 ;
        RECT 4.165 3.230 4.395 3.620 ;
        RECT 5.895 2.115 6.125 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.525 0.300 1.755 0.690 ;
        RECT 4.165 0.300 4.395 0.690 ;
        RECT 5.895 0.300 6.125 1.385 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.547000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.095 0.980 5.490 3.390 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 2.170 4.075 2.400 ;
        RECT 0.610 1.955 0.840 2.170 ;
        RECT 0.375 1.590 0.840 1.955 ;
        RECT 3.845 1.590 4.075 2.170 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 1.595 2.095 1.940 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.420 1.590 3.500 1.940 ;
    END
  END C
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.000 0.435 3.060 ;
        RECT 0.205 2.770 4.865 3.000 ;
        RECT 0.205 2.715 0.435 2.770 ;
        RECT 0.205 1.150 0.435 1.225 ;
        RECT 4.635 1.150 4.865 2.770 ;
        RECT 0.205 0.920 4.865 1.150 ;
        RECT 0.205 0.840 0.435 0.920 ;
  END
END gf180mcu_as_sc_mcu7t3v3__maj3_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__maj3_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__maj3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 1.525 3.230 1.755 3.620 ;
        RECT 4.165 3.230 4.395 3.620 ;
        RECT 5.895 2.115 6.125 3.620 ;
        RECT 7.495 2.145 7.725 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.830 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.525 0.300 1.755 0.690 ;
        RECT 4.165 0.300 4.395 0.690 ;
        RECT 5.895 0.300 6.125 1.385 ;
        RECT 7.495 0.300 7.725 1.410 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.784600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.095 1.885 5.490 3.390 ;
        RECT 6.695 1.885 6.990 3.390 ;
        RECT 5.095 1.655 6.990 1.885 ;
        RECT 5.095 0.980 5.490 1.655 ;
        RECT 6.695 0.980 6.990 1.655 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.610 2.170 4.075 2.400 ;
        RECT 0.610 1.955 0.840 2.170 ;
        RECT 0.375 1.590 0.840 1.955 ;
        RECT 3.845 1.590 4.075 2.170 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.100 1.595 2.095 1.940 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.420 1.590 3.500 1.940 ;
    END
  END C
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.000 0.435 3.060 ;
        RECT 0.205 2.770 4.865 3.000 ;
        RECT 0.205 2.715 0.435 2.770 ;
        RECT 0.205 1.150 0.435 1.225 ;
        RECT 4.635 1.150 4.865 2.770 ;
        RECT 0.205 0.920 4.865 1.150 ;
        RECT 0.205 0.840 0.435 0.920 ;
  END
END gf180mcu_as_sc_mcu7t3v3__maj3_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__mux2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.720 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.720 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 4.425 3.230 4.655 3.620 ;
        RECT 6.045 2.165 6.275 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 7.150 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.150 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 4.425 0.300 4.655 0.690 ;
        RECT 6.045 0.300 6.275 1.415 ;
        RECT 0.000 -0.300 6.720 0.300 ;
    END
  END VSS
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 1.570 1.000 2.240 ;
        RECT 0.705 1.225 0.935 1.570 ;
        RECT 2.105 1.225 2.335 1.940 ;
        RECT 3.360 1.570 3.720 2.540 ;
        RECT 3.425 1.225 3.655 1.570 ;
        RECT 0.705 0.995 3.655 1.225 ;
    END
  END S
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.570 1.800 2.540 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.960 1.570 4.320 2.540 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.285200 ;
    PORT
      LAYER Metal1 ;
        RECT 5.245 0.990 5.575 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.000 0.435 3.390 ;
        RECT 2.720 3.160 3.775 3.390 ;
        RECT 3.545 3.000 3.775 3.160 ;
        RECT 0.205 2.770 2.485 3.000 ;
        RECT 3.545 2.770 5.015 3.000 ;
        RECT 0.205 0.990 0.435 2.770 ;
        RECT 2.255 2.550 2.485 2.770 ;
        RECT 2.255 2.320 2.940 2.550 ;
        RECT 2.710 1.570 2.940 2.320 ;
        RECT 4.785 1.150 5.015 2.770 ;
        RECT 3.965 0.920 5.015 1.150 ;
        RECT 3.965 0.760 4.195 0.920 ;
        RECT 2.205 0.530 4.195 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__mux2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__mux2_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 4.425 3.230 4.655 3.620 ;
        RECT 6.045 2.165 6.275 3.620 ;
        RECT 7.645 2.165 7.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.830 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 4.425 0.300 4.655 0.690 ;
        RECT 6.045 0.300 6.275 1.415 ;
        RECT 7.645 0.300 7.875 1.415 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 1.570 1.000 2.240 ;
        RECT 0.705 1.225 0.935 1.570 ;
        RECT 2.105 1.225 2.335 1.940 ;
        RECT 3.360 1.570 3.720 2.540 ;
        RECT 3.425 1.225 3.655 1.570 ;
        RECT 0.705 0.995 3.655 1.225 ;
    END
  END S
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.570 1.800 2.540 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 3.960 1.570 4.320 2.540 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.522800 ;
    PORT
      LAYER Metal1 ;
        RECT 5.245 1.890 5.575 3.390 ;
        RECT 6.845 1.890 7.175 3.390 ;
        RECT 5.245 1.660 7.175 1.890 ;
        RECT 5.245 0.990 5.575 1.660 ;
        RECT 6.845 0.990 7.175 1.660 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.000 0.435 3.390 ;
        RECT 2.720 3.160 3.775 3.390 ;
        RECT 3.545 3.000 3.775 3.160 ;
        RECT 0.205 2.770 2.485 3.000 ;
        RECT 3.545 2.770 5.015 3.000 ;
        RECT 0.205 0.990 0.435 2.770 ;
        RECT 2.255 2.550 2.485 2.770 ;
        RECT 2.255 2.320 2.940 2.550 ;
        RECT 2.710 1.570 2.940 2.320 ;
        RECT 4.785 1.150 5.015 2.770 ;
        RECT 3.965 0.920 5.015 1.150 ;
        RECT 3.965 0.760 4.195 0.920 ;
        RECT 2.205 0.530 4.195 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__mux2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 0.205 2.840 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.410 3.230 3.640 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.955200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 3.000 1.235 3.160 ;
        RECT 2.605 3.000 2.835 3.160 ;
        RECT 1.005 2.770 3.635 3.000 ;
        RECT 2.605 1.320 2.835 1.330 ;
        RECT 3.165 1.320 3.635 2.770 ;
        RECT 2.605 1.050 3.635 1.320 ;
        RECT 2.605 0.990 2.835 1.050 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.130 1.610 2.935 2.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 1.615 1.660 2.020 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 0.205 0.920 2.035 1.150 ;
        RECT 0.205 0.805 0.435 0.920 ;
        RECT 1.805 0.760 2.035 0.920 ;
        RECT 1.805 0.530 3.690 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand2_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 0.205 2.235 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 3.230 3.635 3.620 ;
        RECT 5.005 3.230 5.235 3.620 ;
        RECT 6.605 2.135 6.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.415 1.770 7.725 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 2.605 0.300 2.835 0.690 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.910400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.805 2.710 6.035 3.390 ;
        RECT 0.820 2.480 6.035 2.710 ;
        RECT 5.805 2.265 6.035 2.480 ;
        RECT 5.805 1.245 6.165 2.265 ;
        RECT 4.085 1.015 6.165 1.245 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 1.600 3.145 2.055 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.895 1.595 5.540 2.050 ;
    END
  END B
  OBS
      LAYER Metal1 ;
        RECT 0.205 1.245 0.435 1.315 ;
        RECT 1.805 1.245 2.035 1.315 ;
        RECT 3.405 1.245 3.635 1.315 ;
        RECT 0.205 1.015 3.635 1.245 ;
        RECT 0.205 0.950 0.435 1.015 ;
        RECT 1.805 0.950 2.035 1.015 ;
        RECT 3.405 0.760 3.635 1.015 ;
        RECT 3.405 0.530 6.890 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand2b_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.445 2.360 0.675 3.620 ;
        RECT 1.885 2.360 2.115 3.620 ;
        RECT 3.485 3.230 3.715 3.620 ;
        RECT 5.090 3.230 5.320 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.300 0.675 1.365 ;
        RECT 2.685 0.300 2.915 0.690 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.955200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.685 3.000 2.915 3.160 ;
        RECT 4.285 3.000 4.515 3.160 ;
        RECT 2.685 2.770 5.315 3.000 ;
        RECT 4.285 1.320 4.515 1.330 ;
        RECT 4.845 1.320 5.315 2.770 ;
        RECT 4.285 1.050 5.315 1.320 ;
        RECT 4.285 0.990 4.515 1.050 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.810 1.610 4.615 2.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.310 1.595 1.010 1.945 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.915 1.475 3.390 ;
        RECT 2.180 1.915 2.480 2.020 ;
        RECT 1.245 1.685 2.480 1.915 ;
        RECT 1.245 0.990 1.475 1.685 ;
        RECT 2.180 1.615 2.480 1.685 ;
        RECT 1.885 0.920 3.715 1.150 ;
        RECT 1.885 0.805 2.115 0.920 ;
        RECT 3.485 0.760 3.715 0.920 ;
        RECT 3.485 0.530 5.370 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand2b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand2b_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 0.445 2.180 0.675 3.620 ;
        RECT 1.885 2.235 2.115 3.620 ;
        RECT 3.485 3.230 3.715 3.620 ;
        RECT 5.085 3.230 5.315 3.620 ;
        RECT 6.685 3.230 6.915 3.620 ;
        RECT 8.285 2.135 8.515 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.300 0.675 1.350 ;
        RECT 2.685 0.300 2.915 0.690 ;
        RECT 4.285 0.300 4.515 0.690 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.910400 ;
    PORT
      LAYER Metal1 ;
        RECT 7.485 2.710 7.715 3.390 ;
        RECT 2.500 2.480 7.715 2.710 ;
        RECT 7.485 2.265 7.715 2.480 ;
        RECT 7.485 1.245 7.845 2.265 ;
        RECT 5.765 1.015 7.845 1.245 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 1.580 1.015 1.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.575 1.595 7.220 2.050 ;
    END
  END B
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.880 1.475 3.390 ;
        RECT 2.260 1.880 2.555 1.930 ;
        RECT 1.245 1.650 2.555 1.880 ;
        RECT 1.245 0.975 1.475 1.650 ;
        RECT 2.260 1.590 2.555 1.650 ;
        RECT 1.885 1.245 2.115 1.315 ;
        RECT 3.485 1.245 3.715 1.315 ;
        RECT 5.085 1.245 5.315 1.315 ;
        RECT 1.885 1.015 5.315 1.245 ;
        RECT 1.885 0.950 2.115 1.015 ;
        RECT 3.485 0.950 3.715 1.015 ;
        RECT 5.085 0.760 5.315 1.015 ;
        RECT 5.085 0.530 8.570 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand2b_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand3_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 0.205 2.300 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 3.230 4.275 3.620 ;
        RECT 5.645 2.210 5.875 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.375 1.585 1.425 1.970 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.975 1.570 3.260 1.955 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.180 1.585 4.580 2.415 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.672800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.580 1.235 3.390 ;
        RECT 2.605 2.875 2.835 3.390 ;
        RECT 4.845 2.875 5.075 3.390 ;
        RECT 2.605 2.750 5.075 2.875 ;
        RECT 2.605 2.645 5.180 2.750 ;
        RECT 2.605 2.580 2.835 2.645 ;
        RECT 1.005 2.350 2.835 2.580 ;
        RECT 4.845 1.255 5.180 2.645 ;
        RECT 4.770 1.025 5.180 1.255 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 1.150 0.435 1.205 ;
        RECT 0.205 0.920 2.035 1.150 ;
        RECT 2.355 0.990 4.275 1.220 ;
        RECT 0.205 0.865 0.435 0.920 ;
        RECT 1.805 0.760 2.035 0.920 ;
        RECT 4.045 0.760 4.275 0.990 ;
        RECT 1.805 0.530 3.690 0.760 ;
        RECT 4.045 0.530 5.930 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand3_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nand4_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
        RECT 0.205 2.300 0.435 3.620 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 3.230 4.275 3.620 ;
        RECT 5.645 3.230 5.875 3.620 ;
        RECT 7.245 2.150 7.475 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.270 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.270 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.375 1.585 1.425 1.970 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.975 1.570 3.260 1.955 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.180 1.585 4.580 2.415 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 5.780 1.585 6.180 2.415 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.390400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.580 1.235 3.390 ;
        RECT 2.605 2.875 2.835 3.390 ;
        RECT 4.845 2.875 5.075 3.045 ;
        RECT 6.445 2.875 6.675 3.045 ;
        RECT 2.605 2.645 6.675 2.875 ;
        RECT 2.605 2.580 2.835 2.645 ;
        RECT 1.005 2.350 2.835 2.580 ;
        RECT 6.445 2.560 6.675 2.645 ;
        RECT 6.445 0.990 6.875 2.560 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 1.150 0.435 1.205 ;
        RECT 0.205 0.920 2.035 1.150 ;
        RECT 2.355 0.990 5.130 1.220 ;
        RECT 0.205 0.865 0.435 0.920 ;
        RECT 1.805 0.760 2.035 0.920 ;
        RECT 1.805 0.530 3.690 0.760 ;
        RECT 3.990 0.530 7.530 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nand4_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nor2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.757600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.545 2.285 3.635 2.555 ;
        RECT 2.605 1.320 2.835 1.330 ;
        RECT 3.165 1.320 3.635 2.285 ;
        RECT 2.605 1.275 3.635 1.320 ;
        RECT 1.005 1.050 3.635 1.275 ;
        RECT 1.005 1.045 2.835 1.050 ;
        RECT 1.005 0.935 1.235 1.045 ;
        RECT 2.605 0.990 2.835 1.045 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.130 1.610 2.935 2.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.500 1.615 1.660 2.020 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.750 3.160 3.690 3.390 ;
        RECT 0.205 2.925 0.435 3.040 ;
        RECT 1.750 2.925 1.980 3.160 ;
        RECT 0.205 2.695 1.980 2.925 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nor2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nor2_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.280 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.280 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 2.605 3.230 2.835 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 7.710 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 7.710 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.370 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 5.005 0.300 5.235 0.690 ;
        RECT 6.605 0.300 6.835 1.370 ;
        RECT 0.000 -0.300 7.280 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.515200 ;
    PORT
      LAYER Metal1 ;
        RECT 5.705 2.750 6.135 2.765 ;
        RECT 3.975 2.520 6.135 2.750 ;
        RECT 5.705 1.210 6.135 2.520 ;
        RECT 0.730 0.980 6.135 1.210 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.580 1.565 3.260 1.995 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 3.855 1.565 5.475 1.985 ;
    END
  END B
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.630 0.435 3.390 ;
        RECT 3.405 3.160 6.890 3.390 ;
        RECT 3.405 2.630 3.635 3.160 ;
        RECT 0.205 2.400 3.690 2.630 ;
        RECT 0.205 2.320 0.435 2.400 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nor2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nor2b_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nor2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 0.445 2.595 0.675 3.620 ;
        RECT 2.685 3.230 2.915 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.300 0.675 1.315 ;
        RECT 1.885 0.300 2.115 0.690 ;
        RECT 3.485 0.300 3.715 0.690 ;
        RECT 5.085 0.300 5.315 0.690 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.757600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.845 2.845 5.315 2.930 ;
        RECT 4.225 2.615 5.315 2.845 ;
        RECT 4.845 1.275 5.315 2.615 ;
        RECT 2.685 1.045 5.315 1.275 ;
        RECT 2.685 0.935 2.915 1.045 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.330 1.610 4.615 2.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 1.975 0.775 2.365 ;
        RECT 0.415 1.545 0.975 1.975 ;
    END
  END A
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.935 1.475 3.390 ;
        RECT 3.430 3.160 5.370 3.390 ;
        RECT 1.885 2.925 2.115 3.040 ;
        RECT 3.430 2.925 3.660 3.160 ;
        RECT 1.885 2.695 3.660 2.925 ;
        RECT 2.180 1.935 2.500 2.020 ;
        RECT 1.245 1.705 2.500 1.935 ;
        RECT 1.245 0.990 1.475 1.705 ;
        RECT 2.180 1.615 2.500 1.705 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nor2b_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nor2b_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nor2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.960 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.960 4.220 ;
        RECT 0.445 2.615 0.675 3.620 ;
        RECT 2.685 3.230 2.915 3.620 ;
        RECT 4.285 3.230 4.515 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 9.390 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 9.390 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 0.300 0.675 1.310 ;
        RECT 1.885 0.300 2.115 1.370 ;
        RECT 3.485 0.300 3.715 0.690 ;
        RECT 5.085 0.300 5.315 0.690 ;
        RECT 6.685 0.300 6.915 0.690 ;
        RECT 8.285 0.300 8.515 1.370 ;
        RECT 0.000 -0.300 8.960 0.300 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.515200 ;
    PORT
      LAYER Metal1 ;
        RECT 7.385 2.750 7.815 2.930 ;
        RECT 5.655 2.520 7.815 2.750 ;
        RECT 7.385 1.210 7.815 2.520 ;
        RECT 2.410 0.980 7.815 1.210 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.410 1.955 0.755 2.385 ;
        RECT 0.410 1.545 0.970 1.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.665600 ;
    PORT
      LAYER Metal1 ;
        RECT 5.535 1.565 7.155 1.985 ;
    END
  END B
  OBS
      LAYER Metal1 ;
        RECT 1.245 1.895 1.475 3.390 ;
        RECT 1.885 2.630 2.115 3.390 ;
        RECT 5.085 3.160 8.570 3.390 ;
        RECT 5.085 2.630 5.315 3.160 ;
        RECT 1.885 2.400 5.370 2.630 ;
        RECT 1.885 2.320 2.115 2.400 ;
        RECT 2.225 1.895 2.550 1.955 ;
        RECT 1.245 1.665 2.550 1.895 ;
        RECT 1.245 0.990 1.475 1.665 ;
        RECT 2.225 1.610 2.550 1.665 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nor2b_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__nor3_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.160 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 6.160 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.590 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.590 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.355 ;
        RECT 1.805 0.300 2.035 0.715 ;
        RECT 3.405 0.300 4.275 0.715 ;
        RECT 5.645 0.300 5.875 1.370 ;
        RECT 0.000 -0.300 6.160 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.375 1.585 1.425 1.970 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.975 1.570 3.260 1.955 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.180 1.585 4.580 2.415 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.277600 ;
    PORT
      LAYER Metal1 ;
        RECT 4.845 1.255 5.180 2.805 ;
        RECT 1.005 1.025 5.180 1.255 ;
        RECT 1.005 0.835 1.235 1.025 ;
        RECT 2.605 0.830 2.835 1.025 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 1.805 3.125 3.690 3.355 ;
        RECT 0.205 2.875 0.435 2.930 ;
        RECT 1.805 2.875 2.035 3.125 ;
        RECT 4.045 3.100 5.875 3.330 ;
        RECT 4.045 2.875 4.275 3.100 ;
        RECT 0.205 2.650 2.035 2.875 ;
        RECT 0.205 2.645 1.910 2.650 ;
        RECT 2.550 2.645 4.275 2.875 ;
        RECT 0.205 2.590 0.435 2.645 ;
        RECT 5.645 2.125 5.875 3.100 ;
  END
END gf180mcu_as_sc_mcu7t3v3__nor3_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__oai211_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__oai211_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.400 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 8.400 4.220 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 4.325 3.230 4.555 3.620 ;
        RECT 5.925 3.230 6.155 3.620 ;
        RECT 7.525 3.230 7.755 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 8.830 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 8.830 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 0.690 ;
        RECT 0.000 -0.300 8.400 0.300 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.620 1.580 1.585 1.985 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 1.565 3.200 1.970 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 4.650 1.985 4.990 2.470 ;
        RECT 4.650 1.585 5.780 1.985 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.672800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.525 2.700 7.050 2.930 ;
        RECT 6.725 0.990 7.050 2.700 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 7.410 1.565 8.140 1.965 ;
    END
  END D
  OBS
      LAYER Metal1 ;
        RECT 0.205 3.000 0.435 3.230 ;
        RECT 1.805 3.160 3.690 3.390 ;
        RECT 1.805 3.000 2.035 3.160 ;
        RECT 0.205 2.770 2.035 3.000 ;
        RECT 4.325 1.220 4.555 1.330 ;
        RECT 0.930 0.925 4.095 1.155 ;
        RECT 4.325 0.990 6.155 1.220 ;
        RECT 3.865 0.760 4.095 0.925 ;
        RECT 5.925 0.760 6.155 0.990 ;
        RECT 3.865 0.530 5.415 0.760 ;
        RECT 5.925 0.530 7.840 0.760 ;
  END
END gf180mcu_as_sc_mcu7t3v3__oai211_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__or2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.920 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.920 4.220 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 2.150 3.635 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 4.350 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 4.350 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 1.450 ;
        RECT 0.000 -0.300 3.920 0.300 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.555 1.660 2.540 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.560 0.860 1.985 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.605 0.920 3.035 3.390 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.770 2.120 3.000 ;
        RECT 0.205 2.640 0.435 2.770 ;
        RECT 1.890 1.980 2.120 2.770 ;
        RECT 1.890 1.555 2.195 1.980 ;
        RECT 1.890 1.150 2.120 1.555 ;
        RECT 0.940 0.920 2.120 1.150 ;
  END
END gf180mcu_as_sc_mcu7t3v3__or2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__or2_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 5.600 4.220 ;
        RECT 1.805 3.230 2.035 3.620 ;
        RECT 3.405 2.150 3.635 3.620 ;
        RECT 5.005 2.150 5.235 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 6.030 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 6.030 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 0.690 ;
        RECT 1.805 0.300 2.035 0.690 ;
        RECT 3.405 0.300 3.635 1.425 ;
        RECT 5.005 0.300 5.235 1.425 ;
        RECT 0.000 -0.300 5.600 0.300 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.555 1.660 2.540 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 1.560 0.860 1.985 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.475200 ;
    PORT
      LAYER Metal1 ;
        RECT 2.605 1.885 2.835 3.390 ;
        RECT 4.205 1.885 4.600 3.390 ;
        RECT 2.605 1.655 4.600 1.885 ;
        RECT 2.605 0.920 2.835 1.655 ;
        RECT 4.205 0.920 4.600 1.655 ;
    END
  END Y
  OBS
      LAYER Metal1 ;
        RECT 0.205 2.770 2.120 3.000 ;
        RECT 0.205 2.640 0.435 2.770 ;
        RECT 1.890 1.980 2.120 2.770 ;
        RECT 1.890 1.555 2.195 1.980 ;
        RECT 1.890 1.150 2.120 1.555 ;
        RECT 0.940 0.920 2.120 1.150 ;
  END
END gf180mcu_as_sc_mcu7t3v3__or2_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__tap_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.120 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 1.550 4.350 ;
      LAYER Metal1 ;
        RECT 0.000 3.620 1.120 4.220 ;
        RECT 0.375 2.235 0.715 3.620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 1.550 1.770 ;
      LAYER Metal1 ;
        RECT 0.375 0.300 0.715 1.380 ;
        RECT 0.000 -0.300 1.120 0.300 ;
    END
  END VSS
END gf180mcu_as_sc_mcu7t3v3__tap_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__tieh_4
  CLASS CORE TIEHIGH ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__tieh_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.205 2.220 0.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.375 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN ONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal1 ;
        RECT 1.005 2.190 1.365 3.390 ;
    END
  END ONE
  OBS
      LAYER Metal1 ;
        RECT 0.570 1.660 1.235 1.895 ;
        RECT 1.005 0.530 1.235 1.660 ;
  END
END gf180mcu_as_sc_mcu7t3v3__tieh_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__tiel_4
  CLASS CORE TIELOW ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__tiel_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
        RECT 0.205 2.220 0.435 3.620 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 1.770 2.670 4.350 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 -0.430 2.670 1.770 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.300 0.435 1.375 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN ZERO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.920 0.530 1.280 1.425 ;
    END
  END ZERO
  OBS
      LAYER Metal1 ;
        RECT 1.005 1.895 1.235 3.390 ;
        RECT 0.570 1.660 1.235 1.895 ;
  END
END gf180mcu_as_sc_mcu7t3v3__tiel_4


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__xnor2_2
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.840 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 7.840 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.920 8.270 4.350 ;
        RECT -0.430 1.770 0.000 3.920 ;
        RECT 0.050 3.670 0.550 3.920 ;
        RECT 7.840 1.770 8.270 3.920 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 0.000 0.000 1.770 ;
        RECT 0.050 0.000 0.550 0.250 ;
        RECT 7.840 0.000 8.270 1.770 ;
        RECT -0.430 -0.430 8.270 0.000 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 7.840 0.300 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.005 1.600 5.440 2.010 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 1.590 1.040 2.655 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.356600 ;
    PORT
      LAYER Metal1 ;
        RECT 6.195 0.990 6.550 3.390 ;
    END
  END Y
  OBS
      LAYER Nwell ;
        RECT 0.000 3.670 0.050 3.920 ;
        RECT 0.550 3.670 7.840 3.920 ;
        RECT 0.000 1.770 7.840 3.670 ;
      LAYER Pwell ;
        RECT 0.000 0.250 7.840 1.770 ;
        RECT 0.000 0.000 0.050 0.250 ;
        RECT 0.550 0.000 7.840 0.250 ;
      LAYER Metal1 ;
        RECT 0.205 3.145 0.435 3.390 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 5.345 3.230 5.575 3.620 ;
        RECT 0.205 2.885 0.755 3.145 ;
        RECT 0.205 1.340 0.435 2.885 ;
        RECT 2.425 2.765 5.965 2.995 ;
        RECT 1.935 2.655 2.195 2.745 ;
        RECT 1.040 2.425 2.195 2.655 ;
        RECT 1.935 2.365 2.195 2.425 ;
        RECT 1.965 1.340 2.195 2.000 ;
        RECT 0.205 1.110 2.195 1.340 ;
        RECT 2.425 1.275 2.655 2.765 ;
        RECT 2.885 2.305 4.775 2.535 ;
        RECT 2.885 1.565 3.115 2.305 ;
        RECT 3.420 1.580 3.715 2.075 ;
        RECT 0.205 0.990 0.435 1.110 ;
        RECT 2.425 1.045 3.210 1.275 ;
        RECT 3.440 1.235 3.700 1.245 ;
        RECT 4.085 1.235 4.315 1.940 ;
        RECT 3.440 1.005 4.315 1.235 ;
        RECT 3.440 0.865 3.700 1.005 ;
        RECT 4.545 0.980 4.775 2.305 ;
        RECT 5.735 1.960 5.965 2.765 ;
        RECT 6.995 2.175 7.225 3.620 ;
        RECT 5.670 1.600 5.965 1.960 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 5.345 0.300 5.575 0.690 ;
        RECT 6.995 0.300 7.225 1.375 ;
      LAYER Metal2 ;
        RECT 0.375 3.155 0.710 3.160 ;
        RECT 1.315 3.155 3.710 3.255 ;
        RECT 0.375 2.975 3.710 3.155 ;
        RECT 0.375 2.875 1.595 2.975 ;
        RECT 0.375 2.870 0.710 2.875 ;
        RECT 1.875 2.365 2.255 2.695 ;
        RECT 1.965 1.190 2.245 2.365 ;
        RECT 3.430 2.030 3.710 2.975 ;
        RECT 3.420 1.695 3.715 2.030 ;
        RECT 3.410 1.190 3.730 1.245 ;
        RECT 1.965 0.910 3.730 1.190 ;
        RECT 3.410 0.865 3.730 0.910 ;
  END
END gf180mcu_as_sc_mcu7t3v3__xnor2_2


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t3v3__xnor2_4
  CLASS CORE ;
  FOREIGN gf180mcu_as_sc_mcu7t3v3__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.520 BY 3.920 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 9.520 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.920 9.950 4.350 ;
        RECT -0.430 1.770 0.000 3.920 ;
        RECT 0.050 3.670 0.550 3.920 ;
        RECT 9.520 1.770 9.950 3.920 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT -0.430 0.000 0.000 1.770 ;
        RECT 0.050 0.000 0.550 0.250 ;
        RECT 9.520 0.000 9.950 1.770 ;
        RECT -0.430 -0.430 9.950 0.000 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 9.520 0.300 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    PORT
      LAYER Metal1 ;
        RECT 5.005 1.600 5.440 2.010 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.332800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.665 1.590 1.040 2.655 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.594200 ;
    PORT
      LAYER Metal1 ;
        RECT 6.195 0.990 6.550 3.390 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 7.795 0.990 8.095 3.390 ;
    END
  END Y
  OBS
      LAYER Nwell ;
        RECT 0.000 3.670 0.050 3.920 ;
        RECT 0.550 3.670 9.520 3.920 ;
        RECT 0.000 1.770 9.520 3.670 ;
      LAYER Pwell ;
        RECT 0.000 0.250 9.520 1.770 ;
        RECT 0.000 0.000 0.050 0.250 ;
        RECT 0.550 0.000 9.520 0.250 ;
      LAYER Metal1 ;
        RECT 0.205 3.145 0.435 3.390 ;
        RECT 1.005 3.230 1.235 3.620 ;
        RECT 5.345 3.230 5.575 3.620 ;
        RECT 0.205 2.885 0.755 3.145 ;
        RECT 0.205 1.340 0.435 2.885 ;
        RECT 2.425 2.765 5.965 2.995 ;
        RECT 1.935 2.655 2.195 2.745 ;
        RECT 1.040 2.425 2.195 2.655 ;
        RECT 1.935 2.365 2.195 2.425 ;
        RECT 1.965 1.340 2.195 2.000 ;
        RECT 0.205 1.110 2.195 1.340 ;
        RECT 2.425 1.275 2.655 2.765 ;
        RECT 2.885 2.305 4.775 2.535 ;
        RECT 2.885 1.565 3.115 2.305 ;
        RECT 3.420 1.580 3.715 2.075 ;
        RECT 0.205 0.990 0.435 1.110 ;
        RECT 2.425 1.045 3.210 1.275 ;
        RECT 3.440 1.235 3.700 1.245 ;
        RECT 4.085 1.235 4.315 1.940 ;
        RECT 3.440 1.005 4.315 1.235 ;
        RECT 3.440 0.865 3.700 1.005 ;
        RECT 4.545 0.980 4.775 2.305 ;
        RECT 5.735 1.960 5.965 2.765 ;
        RECT 6.995 2.175 7.225 3.620 ;
        RECT 8.595 2.170 8.825 3.620 ;
        RECT 5.670 1.600 5.965 1.960 ;
        RECT 6.550 1.665 7.795 1.895 ;
        RECT 1.005 0.300 1.235 0.690 ;
        RECT 5.345 0.300 5.575 0.690 ;
        RECT 6.995 0.300 7.225 1.375 ;
        RECT 8.595 0.300 8.825 1.375 ;
      LAYER Metal2 ;
        RECT 0.375 3.155 0.710 3.160 ;
        RECT 1.315 3.155 3.710 3.255 ;
        RECT 0.375 2.975 3.710 3.155 ;
        RECT 0.375 2.875 1.595 2.975 ;
        RECT 0.375 2.870 0.710 2.875 ;
        RECT 1.875 2.365 2.255 2.695 ;
        RECT 1.965 1.190 2.245 2.365 ;
        RECT 3.430 2.030 3.710 2.975 ;
        RECT 3.420 1.695 3.715 2.030 ;
        RECT 3.410 1.190 3.730 1.245 ;
        RECT 1.965 0.910 3.730 1.190 ;
        RECT 3.410 0.865 3.730 0.910 ;
  END
END gf180mcu_as_sc_mcu7t3v3__xnor2_4


END LIBRARY
