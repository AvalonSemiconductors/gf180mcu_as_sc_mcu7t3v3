magic
tech gf180mcuD
magscale 1 10
timestamp 1753272495
<< nwell >>
rect -86 354 1430 870
<< pwell >>
rect -86 -86 1430 354
<< nmos >>
rect 116 68 172 268
rect 220 68 276 268
rect 380 68 436 268
rect 484 68 540 268
rect 644 68 700 268
rect 748 68 804 268
rect 908 68 964 268
rect 1094 68 1150 268
<< pmos >>
rect 116 440 172 716
rect 220 440 276 716
rect 380 440 436 716
rect 484 440 540 716
rect 644 440 700 716
rect 748 440 804 716
rect 908 440 964 716
rect 1094 440 1150 716
<< ndiff >>
rect 28 230 116 268
rect 28 184 41 230
rect 87 184 116 230
rect 28 68 116 184
rect 172 68 220 268
rect 276 127 380 268
rect 276 81 305 127
rect 351 81 380 127
rect 276 68 380 81
rect 436 68 484 268
rect 540 230 644 268
rect 540 184 569 230
rect 615 184 644 230
rect 540 68 644 184
rect 700 68 748 268
rect 804 127 908 268
rect 804 81 833 127
rect 879 81 908 127
rect 804 68 908 81
rect 964 255 1094 268
rect 964 209 1019 255
rect 1065 209 1094 255
rect 964 68 1094 209
rect 1150 255 1316 268
rect 1150 81 1179 255
rect 1225 81 1316 255
rect 1150 68 1316 81
<< pdiff >>
rect 28 600 116 716
rect 28 554 41 600
rect 87 554 116 600
rect 28 440 116 554
rect 172 440 220 716
rect 276 703 380 716
rect 276 657 305 703
rect 351 657 380 703
rect 276 440 380 657
rect 436 440 484 716
rect 540 600 644 716
rect 540 554 569 600
rect 615 554 644 600
rect 540 440 644 554
rect 700 440 748 716
rect 804 703 908 716
rect 804 657 833 703
rect 879 657 908 703
rect 804 440 908 657
rect 964 667 1094 716
rect 964 453 1019 667
rect 1065 453 1094 667
rect 964 440 1094 453
rect 1150 703 1316 716
rect 1150 453 1179 703
rect 1225 453 1316 703
rect 1150 440 1316 453
<< ndiffc >>
rect 41 184 87 230
rect 305 81 351 127
rect 569 184 615 230
rect 833 81 879 127
rect 1019 209 1065 255
rect 1179 81 1225 255
<< pdiffc >>
rect 41 554 87 600
rect 305 657 351 703
rect 569 554 615 600
rect 833 657 879 703
rect 1019 453 1065 667
rect 1179 453 1225 703
<< polysilicon >>
rect 116 716 172 760
rect 220 716 276 760
rect 380 716 436 760
rect 484 716 540 760
rect 644 716 700 760
rect 748 716 804 760
rect 908 716 964 760
rect 1094 716 1150 760
rect 116 391 172 440
rect 75 377 172 391
rect 75 331 98 377
rect 144 331 172 377
rect 75 318 172 331
rect 116 268 172 318
rect 220 391 276 440
rect 380 391 436 440
rect 220 378 436 391
rect 220 332 233 378
rect 412 332 436 378
rect 220 319 436 332
rect 220 268 276 319
rect 380 268 436 319
rect 484 390 540 440
rect 644 390 700 440
rect 484 377 700 390
rect 484 331 497 377
rect 687 331 700 377
rect 484 318 700 331
rect 484 268 540 318
rect 644 268 700 318
rect 748 391 804 440
rect 748 377 834 391
rect 748 331 769 377
rect 815 331 834 377
rect 748 318 834 331
rect 908 390 964 440
rect 1094 390 1150 440
rect 908 377 1150 390
rect 908 331 927 377
rect 973 331 1150 377
rect 908 318 1150 331
rect 748 268 804 318
rect 908 268 964 318
rect 1094 268 1150 318
rect 116 24 172 68
rect 220 24 276 68
rect 380 24 436 68
rect 484 24 540 68
rect 644 24 700 68
rect 748 24 804 68
rect 908 24 964 68
rect 1094 24 1150 68
<< polycontact >>
rect 98 331 144 377
rect 233 332 412 378
rect 497 331 687 377
rect 769 331 815 377
rect 927 331 973 377
<< metal1 >>
rect 0 724 1344 844
rect 305 703 351 724
rect 305 646 351 657
rect 833 703 879 724
rect 1179 703 1225 724
rect 833 646 879 657
rect 1019 667 1098 678
rect 41 600 87 612
rect 87 554 569 600
rect 615 554 973 600
rect 41 543 87 554
rect 122 434 815 480
rect 122 391 168 434
rect 75 377 168 391
rect 75 331 98 377
rect 144 331 168 377
rect 75 318 168 331
rect 220 378 419 388
rect 220 332 233 378
rect 412 332 419 378
rect 220 319 419 332
rect 484 377 700 388
rect 484 331 497 377
rect 687 331 700 377
rect 484 318 700 331
rect 769 377 815 434
rect 769 318 815 331
rect 927 377 973 554
rect 41 230 87 245
rect 927 230 973 331
rect 87 184 569 230
rect 615 184 973 230
rect 1065 453 1098 667
rect 1019 255 1098 453
rect 1179 423 1225 453
rect 1065 209 1098 255
rect 1019 196 1098 209
rect 1179 255 1225 277
rect 41 168 87 184
rect 305 127 351 138
rect 305 60 351 81
rect 833 127 879 138
rect 833 60 879 81
rect 1179 60 1225 81
rect 0 -60 1344 60
<< labels >>
flabel metal1 s 0 724 1344 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1344 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 1019 196 1098 678 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 75 318 168 391 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 220 319 419 388 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 484 318 700 388 0 FreeSans 200 0 0 0 C
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1344 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1360 354
string MASKHINTS_PPLUS -16 354 1360 830
<< end >>
