magic
tech gf180mcuD
magscale 1 10
timestamp 1752061857
<< nwell >>
rect -86 354 1878 870
<< pwell >>
rect -86 -86 1878 354
<< nmos >>
rect 164 68 220 268
rect 452 68 508 268
rect 612 68 668 268
rect 772 68 828 268
rect 932 68 988 268
rect 1092 68 1148 268
rect 1252 68 1308 268
rect 1412 68 1468 268
rect 1572 68 1628 268
<< pmos >>
rect 164 440 220 716
rect 452 440 508 716
rect 612 440 668 716
rect 772 440 828 716
rect 932 440 988 716
rect 1092 440 1148 716
rect 1252 440 1308 716
rect 1412 440 1468 716
rect 1572 440 1628 716
<< ndiff >>
rect 75 244 164 268
rect 75 81 89 244
rect 135 81 164 244
rect 75 68 164 81
rect 220 255 308 268
rect 220 209 249 255
rect 295 209 308 255
rect 220 68 308 209
rect 364 255 452 268
rect 364 81 377 255
rect 423 81 452 255
rect 364 68 452 81
rect 508 242 612 268
rect 508 196 537 242
rect 583 196 612 242
rect 508 68 612 196
rect 668 127 772 268
rect 668 81 697 127
rect 743 81 772 127
rect 668 68 772 81
rect 828 242 932 268
rect 828 196 857 242
rect 903 196 932 242
rect 828 68 932 196
rect 988 127 1092 268
rect 988 81 1017 127
rect 1063 81 1092 127
rect 988 68 1092 81
rect 1148 242 1252 268
rect 1148 196 1177 242
rect 1223 196 1252 242
rect 1148 68 1252 196
rect 1308 127 1412 268
rect 1308 81 1337 127
rect 1383 81 1412 127
rect 1308 68 1412 81
rect 1468 242 1572 268
rect 1468 196 1497 242
rect 1543 196 1572 242
rect 1468 68 1572 196
rect 1628 255 1764 268
rect 1628 81 1657 255
rect 1703 81 1764 255
rect 1628 68 1764 81
<< pdiff >>
rect 75 703 164 716
rect 75 534 89 703
rect 135 534 164 703
rect 75 440 164 534
rect 220 667 308 716
rect 220 453 249 667
rect 295 453 308 667
rect 220 440 308 453
rect 364 667 452 716
rect 364 480 377 667
rect 423 480 452 667
rect 364 440 452 480
rect 508 703 612 716
rect 508 657 537 703
rect 583 657 612 703
rect 508 440 612 657
rect 668 526 772 716
rect 668 480 697 526
rect 743 480 772 526
rect 668 440 772 480
rect 828 703 932 716
rect 828 657 857 703
rect 903 657 932 703
rect 828 440 932 657
rect 988 667 1092 716
rect 988 480 1017 667
rect 1063 480 1092 667
rect 988 440 1092 480
rect 1148 550 1252 716
rect 1148 504 1177 550
rect 1223 504 1252 550
rect 1148 440 1252 504
rect 1308 678 1412 716
rect 1308 632 1337 678
rect 1383 632 1412 678
rect 1308 440 1412 632
rect 1468 550 1572 716
rect 1468 504 1497 550
rect 1543 504 1572 550
rect 1468 440 1572 504
rect 1628 678 1764 716
rect 1628 632 1657 678
rect 1703 632 1764 678
rect 1628 440 1764 632
<< ndiffc >>
rect 89 81 135 244
rect 249 209 295 255
rect 377 81 423 255
rect 537 196 583 242
rect 697 81 743 127
rect 857 196 903 242
rect 1017 81 1063 127
rect 1177 196 1223 242
rect 1337 81 1383 127
rect 1497 196 1543 242
rect 1657 81 1703 255
<< pdiffc >>
rect 89 534 135 703
rect 249 453 295 667
rect 377 480 423 667
rect 537 657 583 703
rect 697 480 743 526
rect 857 657 903 703
rect 1017 480 1063 667
rect 1177 504 1223 550
rect 1337 632 1383 678
rect 1497 504 1543 550
rect 1657 632 1703 678
<< polysilicon >>
rect 164 716 220 760
rect 452 716 508 760
rect 612 716 668 760
rect 772 716 828 760
rect 932 716 988 760
rect 1092 716 1148 760
rect 1252 716 1308 760
rect 1412 716 1468 760
rect 1572 716 1628 760
rect 164 392 220 440
rect 452 393 508 440
rect 612 393 668 440
rect 772 393 828 440
rect 932 393 988 440
rect 132 379 220 392
rect 132 333 148 379
rect 194 333 220 379
rect 132 320 220 333
rect 445 380 988 393
rect 445 334 458 380
rect 504 347 988 380
rect 504 334 517 347
rect 445 320 517 334
rect 164 268 220 320
rect 452 268 508 320
rect 612 268 668 347
rect 772 268 828 347
rect 932 268 988 347
rect 1092 393 1148 440
rect 1252 393 1308 440
rect 1412 393 1468 440
rect 1572 393 1628 440
rect 1092 379 1630 393
rect 1092 333 1107 379
rect 1431 333 1630 379
rect 1092 317 1630 333
rect 1092 268 1148 317
rect 1252 268 1308 317
rect 1412 268 1468 317
rect 1572 268 1628 317
rect 164 24 220 68
rect 452 24 508 68
rect 612 24 668 68
rect 772 24 828 68
rect 932 24 988 68
rect 1092 24 1148 68
rect 1252 24 1308 68
rect 1412 24 1468 68
rect 1572 24 1628 68
<< polycontact >>
rect 148 333 194 379
rect 458 334 504 380
rect 1107 333 1431 379
<< metal1 >>
rect 0 724 1792 844
rect 89 703 135 724
rect 537 703 583 724
rect 89 523 135 534
rect 249 667 295 678
rect 82 391 151 477
rect 377 667 423 678
rect 537 646 583 657
rect 857 703 903 724
rect 857 646 903 657
rect 1017 667 1337 678
rect 423 480 697 526
rect 743 480 1017 526
rect 1063 632 1337 667
rect 1383 632 1657 678
rect 1703 632 1714 678
rect 1477 550 1563 586
rect 1063 480 1074 526
rect 1131 504 1177 550
rect 1223 504 1497 550
rect 1543 504 1563 550
rect 377 464 423 480
rect 82 379 194 391
rect 82 333 148 379
rect 82 309 194 333
rect 249 379 295 453
rect 445 380 510 391
rect 445 379 458 380
rect 249 334 458 379
rect 504 334 510 380
rect 249 333 510 334
rect 89 244 135 262
rect 249 255 295 333
rect 445 322 510 333
rect 1107 379 1431 397
rect 1107 313 1431 333
rect 249 198 295 209
rect 377 255 423 274
rect 89 60 135 81
rect 1477 242 1563 504
rect 482 196 537 242
rect 583 196 857 242
rect 903 196 1177 242
rect 1223 196 1497 242
rect 1543 196 1563 242
rect 1657 255 1703 274
rect 377 60 423 81
rect 697 127 743 138
rect 697 60 743 81
rect 1017 127 1063 138
rect 1017 60 1063 81
rect 1337 127 1383 138
rect 1337 60 1383 81
rect 1657 60 1703 81
rect 0 -60 1792 60
<< labels >>
flabel metal1 s 0 724 1792 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1792 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 1477 196 1563 586 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 1107 313 1431 397 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 82 309 194 391 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 82 391 151 477 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1792 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 1878 354
string MASKHINTS_PPLUS -86 354 1878 870
<< end >>
