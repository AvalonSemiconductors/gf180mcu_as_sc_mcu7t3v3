magic
tech gf180mcuD
magscale 1 10
timestamp 1752051650
<< nwell >>
rect -86 354 1878 870
<< pwell >>
rect -86 -86 1878 354
<< nmos >>
rect 164 68 220 268
rect 452 68 508 268
rect 612 68 668 268
rect 772 68 828 268
rect 932 68 988 268
rect 1092 68 1148 268
rect 1252 68 1308 268
rect 1412 68 1468 268
rect 1572 68 1628 268
<< pmos >>
rect 164 440 220 716
rect 452 440 508 716
rect 612 440 668 716
rect 772 440 828 716
rect 932 440 988 716
rect 1092 440 1148 716
rect 1252 440 1308 716
rect 1412 440 1468 716
rect 1572 440 1628 716
<< ndiff >>
rect 76 255 164 268
rect 76 81 89 255
rect 135 81 164 255
rect 76 68 164 81
rect 220 252 308 268
rect 220 206 249 252
rect 295 206 308 252
rect 220 68 308 206
rect 364 249 452 268
rect 364 203 377 249
rect 423 203 452 249
rect 364 68 452 203
rect 508 127 612 268
rect 508 81 537 127
rect 583 81 612 127
rect 508 68 612 81
rect 668 249 772 268
rect 668 203 697 249
rect 743 203 772 249
rect 668 68 772 203
rect 828 127 932 268
rect 828 81 857 127
rect 903 81 932 127
rect 828 68 932 81
rect 988 249 1092 268
rect 988 203 1017 249
rect 1063 203 1092 249
rect 988 68 1092 203
rect 1148 249 1252 268
rect 1148 203 1177 249
rect 1223 203 1252 249
rect 1148 68 1252 203
rect 1308 152 1412 268
rect 1308 106 1337 152
rect 1383 106 1412 152
rect 1308 68 1412 106
rect 1468 249 1572 268
rect 1468 203 1497 249
rect 1543 203 1572 249
rect 1468 68 1572 203
rect 1628 152 1764 268
rect 1628 106 1657 152
rect 1703 106 1764 152
rect 1628 68 1764 106
<< pdiff >>
rect 76 703 164 716
rect 76 453 89 703
rect 135 453 164 703
rect 76 440 164 453
rect 220 667 308 716
rect 220 453 249 667
rect 295 453 308 667
rect 220 440 308 453
rect 364 703 452 716
rect 364 458 377 703
rect 423 458 452 703
rect 364 440 452 458
rect 508 542 612 716
rect 508 496 537 542
rect 583 496 612 542
rect 508 440 612 496
rect 668 703 772 716
rect 668 657 697 703
rect 743 657 772 703
rect 668 440 772 657
rect 828 542 932 716
rect 828 496 857 542
rect 903 496 932 542
rect 828 440 932 496
rect 988 703 1092 716
rect 988 657 1017 703
rect 1063 657 1092 703
rect 988 440 1092 657
rect 1148 542 1252 716
rect 1148 496 1177 542
rect 1223 496 1252 542
rect 1148 440 1252 496
rect 1308 703 1412 716
rect 1308 657 1337 703
rect 1383 657 1412 703
rect 1308 440 1412 657
rect 1468 667 1572 716
rect 1468 453 1497 667
rect 1543 453 1572 667
rect 1468 440 1572 453
rect 1628 703 1764 716
rect 1628 453 1657 703
rect 1703 453 1764 703
rect 1628 440 1764 453
<< ndiffc >>
rect 89 81 135 255
rect 249 206 295 252
rect 377 203 423 249
rect 537 81 583 127
rect 697 203 743 249
rect 857 81 903 127
rect 1017 203 1063 249
rect 1177 203 1223 249
rect 1337 106 1383 152
rect 1497 203 1543 249
rect 1657 106 1703 152
<< pdiffc >>
rect 89 453 135 703
rect 249 453 295 667
rect 377 458 423 703
rect 537 496 583 542
rect 697 657 743 703
rect 857 496 903 542
rect 1017 657 1063 703
rect 1177 496 1223 542
rect 1337 657 1383 703
rect 1497 453 1543 667
rect 1657 453 1703 703
<< polysilicon >>
rect 164 716 220 760
rect 452 716 508 760
rect 612 716 668 760
rect 772 716 828 760
rect 932 716 988 760
rect 1092 716 1148 760
rect 1252 716 1308 760
rect 1412 716 1468 760
rect 1572 716 1628 760
rect 164 390 220 440
rect 131 375 220 390
rect 131 329 146 375
rect 192 329 220 375
rect 131 316 220 329
rect 164 268 220 316
rect 452 389 508 440
rect 452 375 541 389
rect 452 329 465 375
rect 511 372 541 375
rect 612 372 668 440
rect 772 372 828 440
rect 932 372 988 440
rect 511 329 988 372
rect 452 320 988 329
rect 452 315 541 320
rect 452 268 508 315
rect 612 268 668 320
rect 772 268 828 320
rect 932 268 988 320
rect 1092 410 1148 440
rect 1252 410 1308 440
rect 1412 410 1468 440
rect 1572 410 1628 440
rect 1092 391 1628 410
rect 1092 345 1115 391
rect 1444 345 1628 391
rect 1092 319 1628 345
rect 1092 268 1148 319
rect 1252 268 1308 319
rect 1412 268 1468 319
rect 1572 268 1628 319
rect 164 24 220 68
rect 452 24 508 68
rect 612 24 668 68
rect 772 24 828 68
rect 932 24 988 68
rect 1092 24 1148 68
rect 1252 24 1308 68
rect 1412 24 1468 68
rect 1572 24 1628 68
<< polycontact >>
rect 146 329 192 375
rect 465 329 511 375
rect 1115 345 1444 391
<< metal1 >>
rect 0 724 1792 844
rect 89 703 135 724
rect 377 703 423 724
rect 89 436 135 453
rect 249 667 295 678
rect 74 375 203 390
rect 74 329 146 375
rect 192 329 203 375
rect 74 316 203 329
rect 249 376 295 453
rect 697 703 743 724
rect 697 646 743 657
rect 1017 703 1063 724
rect 1017 646 1063 657
rect 1337 703 1383 724
rect 1657 703 1703 724
rect 1337 646 1383 657
rect 1497 667 1543 678
rect 500 496 537 542
rect 583 496 857 542
rect 903 496 1177 542
rect 1223 496 1497 542
rect 377 447 423 458
rect 1115 391 1444 410
rect 452 376 511 386
rect 249 375 511 376
rect 249 330 465 375
rect 89 255 135 270
rect 249 252 295 330
rect 452 329 465 330
rect 452 318 511 329
rect 1115 319 1444 345
rect 249 195 295 206
rect 377 249 423 263
rect 697 249 743 263
rect 1017 249 1063 263
rect 1497 249 1569 453
rect 1657 427 1703 453
rect 423 203 697 249
rect 743 203 1017 249
rect 1153 203 1177 249
rect 1223 203 1497 249
rect 1543 203 1569 249
rect 377 190 423 203
rect 697 190 743 203
rect 1017 152 1063 203
rect 89 60 135 81
rect 537 127 583 138
rect 537 60 583 81
rect 857 127 903 138
rect 1017 106 1337 152
rect 1383 106 1657 152
rect 1703 106 1714 152
rect 857 60 903 81
rect 0 -60 1792 60
<< labels >>
flabel metal1 s 0 724 1792 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1792 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel nwell s 13 734 113 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel metal1 1497 203 1569 453 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 1115 319 1444 410 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 74 316 203 390 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1792 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1808 354
string MASKHINTS_PPLUS -16 354 1808 830
<< end >>
