magic
tech gf180mcuD
magscale 1 10
timestamp 1759934137
<< nwell >>
rect -86 354 1654 870
<< pwell >>
rect -86 -86 1654 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 884 68 940 268
rect 1044 68 1100 268
rect 1204 68 1260 268
rect 1364 68 1420 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 884 440 940 716
rect 1044 440 1100 716
rect 1204 440 1260 716
rect 1364 440 1420 716
<< ndiff >>
rect 28 217 116 268
rect 28 171 41 217
rect 87 171 116 217
rect 28 68 116 171
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 181 436 268
rect 332 135 361 181
rect 407 135 436 181
rect 332 68 436 135
rect 492 255 596 268
rect 492 209 521 255
rect 567 209 596 255
rect 492 68 596 209
rect 652 152 740 268
rect 652 106 681 152
rect 727 106 740 152
rect 652 68 740 106
rect 796 127 884 268
rect 796 81 809 127
rect 855 81 884 127
rect 796 68 884 81
rect 940 163 1044 268
rect 940 117 969 163
rect 1015 117 1044 163
rect 940 68 1044 117
rect 1100 127 1204 268
rect 1100 81 1129 127
rect 1175 81 1204 127
rect 1100 68 1204 81
rect 1260 163 1364 268
rect 1260 117 1289 163
rect 1335 117 1364 163
rect 1260 68 1364 117
rect 1420 127 1513 268
rect 1420 81 1449 127
rect 1495 81 1513 127
rect 1420 68 1513 81
<< pdiff >>
rect 28 703 116 716
rect 28 478 41 703
rect 87 478 116 703
rect 28 440 116 478
rect 172 537 276 716
rect 172 491 201 537
rect 247 491 276 537
rect 172 440 276 491
rect 332 703 436 716
rect 332 657 361 703
rect 407 657 436 703
rect 332 440 436 657
rect 492 548 596 716
rect 492 502 521 548
rect 567 502 596 548
rect 492 440 596 502
rect 652 703 740 716
rect 652 657 681 703
rect 727 657 740 703
rect 652 440 740 657
rect 796 678 884 716
rect 796 632 809 678
rect 855 632 884 678
rect 796 440 884 632
rect 940 570 1044 716
rect 940 524 969 570
rect 1015 524 1044 570
rect 940 440 1044 524
rect 1100 678 1204 716
rect 1100 632 1129 678
rect 1175 632 1204 678
rect 1100 440 1204 632
rect 1260 572 1364 716
rect 1260 526 1289 572
rect 1335 526 1364 572
rect 1260 440 1364 526
rect 1420 678 1513 716
rect 1420 632 1449 678
rect 1495 632 1513 678
rect 1420 440 1513 632
<< ndiffc >>
rect 41 171 87 217
rect 201 81 247 127
rect 361 135 407 181
rect 521 209 567 255
rect 681 106 727 152
rect 809 81 855 127
rect 969 117 1015 163
rect 1129 81 1175 127
rect 1289 117 1335 163
rect 1449 81 1495 127
<< pdiffc >>
rect 41 478 87 703
rect 201 491 247 537
rect 361 657 407 703
rect 521 502 567 548
rect 681 657 727 703
rect 809 632 855 678
rect 969 524 1015 570
rect 1129 632 1175 678
rect 1289 526 1335 572
rect 1449 632 1495 678
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 884 716 940 760
rect 1044 716 1100 760
rect 1204 716 1260 760
rect 1364 716 1420 760
rect 116 413 172 440
rect 75 386 172 413
rect 75 340 99 386
rect 145 385 172 386
rect 276 385 332 440
rect 436 405 492 440
rect 596 405 652 440
rect 145 340 332 385
rect 75 314 332 340
rect 427 384 652 405
rect 884 390 940 440
rect 1044 390 1100 440
rect 427 338 440 384
rect 639 338 652 384
rect 427 319 652 338
rect 116 268 172 314
rect 276 268 332 314
rect 436 268 492 319
rect 596 268 652 319
rect 853 377 1100 390
rect 853 331 866 377
rect 1048 331 1100 377
rect 853 318 1100 331
rect 884 268 940 318
rect 1044 268 1100 318
rect 1204 384 1260 440
rect 1364 408 1420 440
rect 1364 384 1479 408
rect 1204 380 1479 384
rect 1204 334 1389 380
rect 1435 334 1479 380
rect 1204 332 1479 334
rect 1204 268 1260 332
rect 1364 313 1479 332
rect 1364 268 1420 313
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 884 24 940 68
rect 1044 24 1100 68
rect 1204 24 1260 68
rect 1364 24 1420 68
<< polycontact >>
rect 99 340 145 386
rect 440 338 639 384
rect 866 331 1048 377
rect 1389 334 1435 380
<< metal1 >>
rect 0 724 1568 844
rect 41 703 87 724
rect 361 703 407 724
rect 361 646 407 657
rect 681 703 727 724
rect 681 646 727 657
rect 798 632 809 678
rect 855 632 1129 678
rect 1175 632 1449 678
rect 1495 632 1506 678
rect 521 548 969 570
rect 190 491 201 537
rect 247 502 521 537
rect 567 524 969 548
rect 1015 524 1026 570
rect 1147 526 1289 572
rect 1335 526 1346 572
rect 247 491 567 502
rect 41 467 87 478
rect 55 386 171 413
rect 55 340 99 386
rect 145 340 171 386
rect 55 314 171 340
rect 427 384 643 405
rect 427 338 440 384
rect 639 338 643 384
rect 427 319 643 338
rect 853 377 1048 389
rect 853 331 866 377
rect 853 319 1048 331
rect 521 265 567 269
rect 1147 265 1232 526
rect 1364 380 1494 408
rect 1364 334 1389 380
rect 1435 334 1494 380
rect 1364 313 1494 334
rect 521 255 1335 265
rect 41 217 407 239
rect 87 193 407 217
rect 567 219 1335 255
rect 521 198 567 209
rect 41 155 87 171
rect 361 181 407 193
rect 201 127 247 138
rect 969 163 1015 219
rect 407 135 681 152
rect 361 106 681 135
rect 727 106 738 152
rect 809 127 855 138
rect 201 60 247 81
rect 1289 163 1335 219
rect 969 106 1015 117
rect 1129 127 1175 138
rect 809 60 855 81
rect 1289 106 1335 117
rect 1449 127 1495 138
rect 1129 60 1175 81
rect 1449 60 1495 81
rect 0 -60 1568 60
<< labels >>
flabel metal1 s 0 724 1568 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1568 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 55 314 171 413 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 427 319 643 405 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 853 319 1048 389 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 1147 220 1232 572 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel metal1 1364 313 1494 408 0 FreeSans 200 0 0 0 D
port 9 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1584 354
string MASKHINTS_PPLUS -16 354 1584 830
<< end >>
