magic
tech gf180mcuD
magscale 1 10
timestamp 1764158546
<< nwell >>
rect -86 354 1318 870
<< pwell >>
rect -86 -86 1318 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 884 68 940 268
rect 1044 68 1100 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 884 440 940 716
rect 1044 440 1100 716
<< ndiff >>
rect 28 128 116 268
rect 28 82 41 128
rect 87 82 116 128
rect 28 68 116 82
rect 172 68 276 268
rect 332 213 436 268
rect 332 167 361 213
rect 407 167 436 213
rect 332 68 436 167
rect 492 131 596 268
rect 492 85 521 131
rect 567 85 596 131
rect 492 68 596 85
rect 652 220 740 268
rect 652 174 681 220
rect 727 174 740 220
rect 652 68 740 174
rect 796 127 884 268
rect 796 81 809 127
rect 855 81 884 127
rect 796 68 884 81
rect 940 241 1044 268
rect 940 195 969 241
rect 1015 195 1044 241
rect 940 68 1044 195
rect 1100 127 1204 268
rect 1100 81 1129 127
rect 1175 81 1204 127
rect 1100 68 1204 81
<< pdiff >>
rect 28 610 116 716
rect 28 564 41 610
rect 87 564 116 610
rect 28 440 116 564
rect 172 695 276 716
rect 172 649 201 695
rect 247 649 276 695
rect 172 440 276 649
rect 332 610 436 716
rect 332 564 361 610
rect 407 564 436 610
rect 332 440 436 564
rect 492 440 596 716
rect 652 667 740 716
rect 652 515 681 667
rect 727 515 740 667
rect 652 440 740 515
rect 796 698 884 716
rect 796 463 809 698
rect 855 463 884 698
rect 796 440 884 463
rect 940 667 1044 716
rect 940 453 969 667
rect 1015 453 1044 667
rect 940 440 1044 453
rect 1100 695 1204 716
rect 1100 503 1129 695
rect 1175 503 1204 695
rect 1100 440 1204 503
<< ndiffc >>
rect 41 82 87 128
rect 361 167 407 213
rect 521 85 567 131
rect 681 174 727 220
rect 809 81 855 127
rect 969 195 1015 241
rect 1129 81 1175 127
<< pdiffc >>
rect 41 564 87 610
rect 201 649 247 695
rect 361 564 407 610
rect 681 515 727 667
rect 809 463 855 698
rect 969 453 1015 667
rect 1129 503 1175 695
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 884 716 940 760
rect 1044 716 1100 760
rect 116 396 172 440
rect 276 398 332 440
rect 436 399 492 440
rect 596 404 652 440
rect 66 377 172 396
rect 66 331 80 377
rect 126 331 172 377
rect 66 310 172 331
rect 246 377 332 398
rect 246 331 264 377
rect 310 331 332 377
rect 246 313 332 331
rect 406 378 492 399
rect 406 332 421 378
rect 467 332 492 378
rect 406 314 492 332
rect 566 382 652 404
rect 884 391 940 440
rect 1044 391 1100 440
rect 566 336 579 382
rect 625 336 652 382
rect 566 319 652 336
rect 116 268 172 310
rect 276 268 332 313
rect 436 268 492 314
rect 596 268 652 319
rect 825 376 1100 391
rect 825 330 838 376
rect 884 330 1100 376
rect 825 315 1100 330
rect 884 268 940 315
rect 1044 268 1100 315
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 884 24 940 68
rect 1044 24 1100 68
<< polycontact >>
rect 80 331 126 377
rect 264 331 310 377
rect 421 332 467 378
rect 579 336 625 382
rect 838 330 884 376
<< metal1 >>
rect 0 724 1232 844
rect 201 695 247 724
rect 809 698 855 724
rect 201 638 247 649
rect 681 667 727 678
rect 41 610 87 635
rect 361 610 407 632
rect 87 564 361 592
rect 41 546 407 564
rect 727 515 740 550
rect 681 504 740 515
rect 66 377 143 453
rect 66 331 80 377
rect 126 331 143 377
rect 66 310 143 331
rect 246 377 323 451
rect 246 331 264 377
rect 310 331 323 377
rect 246 264 323 331
rect 406 378 483 452
rect 406 332 421 378
rect 467 332 483 378
rect 406 314 483 332
rect 566 382 643 458
rect 566 336 579 382
rect 625 336 643 382
rect 566 307 643 336
rect 694 391 740 504
rect 1129 695 1175 724
rect 809 452 855 463
rect 963 667 1025 678
rect 963 453 969 667
rect 1015 453 1025 667
rect 1129 492 1175 503
rect 694 376 888 391
rect 694 330 838 376
rect 884 330 888 376
rect 694 315 888 330
rect 41 128 87 146
rect 246 119 315 264
rect 694 238 740 315
rect 361 220 740 238
rect 361 213 681 220
rect 407 192 681 213
rect 361 147 407 167
rect 727 174 740 220
rect 681 158 740 174
rect 963 241 1025 453
rect 963 195 969 241
rect 1015 195 1025 241
rect 963 168 1025 195
rect 521 131 567 146
rect 41 60 87 82
rect 521 60 567 85
rect 809 127 855 146
rect 809 60 855 81
rect 1129 127 1175 146
rect 1129 60 1175 81
rect 0 -60 1232 60
<< labels >>
flabel metal1 s 0 724 1232 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1232 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 66 310 143 453 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 246 264 323 451 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 406 314 483 452 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 566 307 643 458 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel metal1 963 168 1025 678 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1232 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1248 354
string MASKHINTS_PPLUS -16 354 1248 830
<< end >>
