magic
tech gf180mcuD
magscale 1 10
timestamp 1751895231
<< nwell >>
rect -86 354 1206 870
<< pwell >>
rect -86 -86 1206 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
<< ndiff >>
rect 28 230 116 268
rect 28 184 41 230
rect 87 184 116 230
rect 28 68 116 184
rect 172 68 276 268
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 251 596 268
rect 492 205 521 251
rect 567 205 596 251
rect 492 68 596 205
rect 652 255 756 268
rect 652 81 681 255
rect 727 81 756 255
rect 652 68 756 81
rect 812 246 916 268
rect 812 200 841 246
rect 887 200 916 246
rect 812 68 916 200
rect 972 255 1092 268
rect 972 81 1001 255
rect 1047 81 1092 255
rect 972 68 1092 81
<< pdiff >>
rect 28 703 116 716
rect 28 657 41 703
rect 87 657 116 703
rect 28 440 116 657
rect 172 600 276 716
rect 172 554 201 600
rect 247 554 276 600
rect 172 440 276 554
rect 332 703 436 716
rect 332 657 361 703
rect 407 657 436 703
rect 332 440 436 657
rect 492 667 596 716
rect 492 453 521 667
rect 567 453 596 667
rect 492 440 596 453
rect 652 703 756 716
rect 652 453 681 703
rect 727 453 756 703
rect 652 440 756 453
rect 812 667 916 716
rect 812 453 841 667
rect 887 453 916 667
rect 812 440 916 453
rect 972 703 1092 716
rect 972 453 1001 703
rect 1047 453 1092 703
rect 972 440 1092 453
<< ndiffc >>
rect 41 184 87 230
rect 361 81 407 127
rect 521 205 567 251
rect 681 81 727 255
rect 841 200 887 246
rect 1001 81 1047 255
<< pdiffc >>
rect 41 657 87 703
rect 201 554 247 600
rect 361 657 407 703
rect 521 453 567 667
rect 681 453 727 703
rect 841 453 887 667
rect 1001 453 1047 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 116 397 172 440
rect 91 379 172 397
rect 276 396 332 440
rect 436 396 492 440
rect 91 333 104 379
rect 150 333 172 379
rect 91 312 172 333
rect 116 268 172 312
rect 251 377 332 396
rect 251 331 271 377
rect 317 331 332 377
rect 251 311 332 331
rect 380 377 492 396
rect 380 331 393 377
rect 439 373 492 377
rect 596 373 652 440
rect 756 373 812 440
rect 916 373 972 440
rect 439 331 972 373
rect 380 330 972 331
rect 380 311 492 330
rect 276 268 332 311
rect 436 268 492 311
rect 596 268 652 330
rect 756 268 812 330
rect 916 268 972 330
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
<< polycontact >>
rect 104 333 150 379
rect 271 331 317 377
rect 393 331 439 377
<< metal1 >>
rect 0 724 1120 844
rect 41 703 87 724
rect 41 646 87 657
rect 361 703 407 724
rect 681 703 727 724
rect 361 646 407 657
rect 521 667 567 678
rect 190 554 201 600
rect 247 554 424 600
rect 41 379 172 397
rect 41 333 104 379
rect 150 333 172 379
rect 41 312 172 333
rect 251 377 332 508
rect 251 331 271 377
rect 317 331 332 377
rect 251 311 332 331
rect 378 396 424 554
rect 378 377 439 396
rect 378 331 393 377
rect 378 311 439 331
rect 521 384 567 453
rect 1001 703 1047 724
rect 681 430 727 453
rect 841 667 920 678
rect 887 453 920 667
rect 841 384 920 453
rect 1001 430 1047 453
rect 521 338 920 384
rect 41 230 87 248
rect 378 230 424 311
rect 87 184 424 230
rect 521 251 567 338
rect 521 184 567 205
rect 681 255 727 290
rect 41 172 87 184
rect 361 127 407 138
rect 361 60 407 81
rect 841 246 920 338
rect 887 200 920 246
rect 841 184 920 200
rect 1001 255 1047 290
rect 681 60 727 81
rect 1001 60 1047 81
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 0 724 1120 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1120 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 251 311 332 508 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel metal1 41 312 172 397 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 841 184 920 678 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1136 354
string MASKHINTS_PPLUS -16 354 1136 830
<< end >>
