magic
tech gf180mcuD
magscale 1 10
timestamp 1752063767
<< nwell >>
rect -86 354 2102 870
<< pwell >>
rect -86 -86 2102 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
rect 1396 68 1452 268
rect 1556 68 1612 268
rect 1716 68 1772 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1396 440 1452 716
rect 1556 440 1612 716
rect 1716 440 1772 716
<< ndiff >>
rect 28 132 116 268
rect 28 86 41 132
rect 87 86 116 132
rect 28 68 116 86
rect 172 255 276 268
rect 172 209 201 255
rect 247 209 276 255
rect 172 68 276 209
rect 332 244 436 268
rect 332 83 361 244
rect 407 83 436 244
rect 332 68 436 83
rect 492 255 596 268
rect 492 209 521 255
rect 567 209 596 255
rect 492 68 596 209
rect 652 255 756 268
rect 652 81 681 255
rect 727 81 756 255
rect 652 68 756 81
rect 812 255 916 268
rect 812 209 841 255
rect 887 209 916 255
rect 812 68 916 209
rect 972 255 1076 268
rect 972 81 1001 255
rect 1047 81 1076 255
rect 972 68 1076 81
rect 1132 255 1236 268
rect 1132 209 1161 255
rect 1207 209 1236 255
rect 1132 68 1236 209
rect 1292 255 1396 268
rect 1292 81 1321 255
rect 1367 81 1396 255
rect 1292 68 1396 81
rect 1452 255 1556 268
rect 1452 209 1481 255
rect 1527 209 1556 255
rect 1452 68 1556 209
rect 1612 254 1716 268
rect 1612 81 1641 254
rect 1687 81 1716 254
rect 1612 68 1716 81
rect 1772 255 1988 268
rect 1772 209 1801 255
rect 1847 209 1988 255
rect 1772 68 1988 209
<< pdiff >>
rect 28 694 116 716
rect 28 648 41 694
rect 87 648 116 694
rect 28 440 116 648
rect 172 667 276 716
rect 172 453 201 667
rect 247 453 276 667
rect 172 440 276 453
rect 332 694 436 716
rect 332 464 361 694
rect 407 464 436 694
rect 332 440 436 464
rect 492 667 596 716
rect 492 453 521 667
rect 567 453 596 667
rect 492 440 596 453
rect 652 696 756 716
rect 652 453 681 696
rect 727 453 756 696
rect 652 440 756 453
rect 812 667 916 716
rect 812 453 841 667
rect 887 453 916 667
rect 812 440 916 453
rect 972 703 1076 716
rect 972 453 1001 703
rect 1047 453 1076 703
rect 972 440 1076 453
rect 1132 667 1236 716
rect 1132 453 1161 667
rect 1207 453 1236 667
rect 1132 440 1236 453
rect 1292 703 1396 716
rect 1292 453 1321 703
rect 1367 453 1396 703
rect 1292 440 1396 453
rect 1452 667 1556 716
rect 1452 453 1481 667
rect 1527 453 1556 667
rect 1452 440 1556 453
rect 1612 703 1716 716
rect 1612 453 1641 703
rect 1687 453 1716 703
rect 1612 440 1716 453
rect 1772 667 1988 716
rect 1772 453 1801 667
rect 1847 453 1988 667
rect 1772 440 1988 453
<< ndiffc >>
rect 41 86 87 132
rect 201 209 247 255
rect 361 83 407 244
rect 521 209 567 255
rect 681 81 727 255
rect 841 209 887 255
rect 1001 81 1047 255
rect 1161 209 1207 255
rect 1321 81 1367 255
rect 1481 209 1527 255
rect 1641 81 1687 254
rect 1801 209 1847 255
<< pdiffc >>
rect 41 648 87 694
rect 201 453 247 667
rect 361 464 407 694
rect 521 453 567 667
rect 681 453 727 696
rect 841 453 887 667
rect 1001 453 1047 703
rect 1161 453 1207 667
rect 1321 453 1367 703
rect 1481 453 1527 667
rect 1641 453 1687 703
rect 1801 453 1847 667
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1396 716 1452 760
rect 1556 716 1612 760
rect 1716 716 1772 760
rect 116 412 172 440
rect 276 412 332 440
rect 74 393 332 412
rect 436 393 492 440
rect 596 399 652 440
rect 756 399 812 440
rect 74 389 492 393
rect 74 343 95 389
rect 141 345 492 389
rect 141 343 332 345
rect 74 322 332 343
rect 116 268 172 322
rect 276 268 332 322
rect 436 268 492 345
rect 544 382 812 399
rect 544 336 557 382
rect 784 378 812 382
rect 916 378 972 440
rect 1076 378 1132 440
rect 1236 378 1292 440
rect 1396 378 1452 440
rect 1556 378 1612 440
rect 1716 378 1772 440
rect 784 336 1772 378
rect 544 332 1772 336
rect 544 322 812 332
rect 596 268 652 322
rect 756 268 812 322
rect 916 268 972 332
rect 1076 268 1132 332
rect 1236 268 1292 332
rect 1396 268 1452 332
rect 1556 268 1612 332
rect 1716 268 1772 332
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1396 24 1452 68
rect 1556 24 1612 68
rect 1716 24 1772 68
<< polycontact >>
rect 95 343 141 389
rect 557 336 784 382
<< metal1 >>
rect 0 724 2016 844
rect 41 694 87 724
rect 361 694 407 724
rect 41 637 87 648
rect 201 667 247 678
rect 41 412 117 481
rect 681 696 727 724
rect 361 453 407 464
rect 521 667 567 678
rect 41 389 154 412
rect 41 343 95 389
rect 141 343 154 389
rect 41 322 154 343
rect 201 407 247 453
rect 521 407 567 453
rect 1001 703 1047 724
rect 681 436 727 453
rect 841 667 887 678
rect 201 399 567 407
rect 201 387 613 399
rect 841 396 887 453
rect 1321 703 1367 724
rect 1001 442 1047 453
rect 1161 667 1207 678
rect 1161 396 1207 453
rect 1641 703 1687 724
rect 1321 442 1367 453
rect 1481 667 1527 678
rect 1481 396 1527 453
rect 1641 442 1687 453
rect 1801 667 1847 678
rect 1801 396 1847 453
rect 201 382 795 387
rect 201 361 557 382
rect 41 291 117 322
rect 201 255 247 361
rect 521 336 557 361
rect 784 336 795 382
rect 521 332 795 336
rect 521 322 613 332
rect 521 255 567 322
rect 841 314 1847 396
rect 201 198 247 209
rect 361 244 407 255
rect 41 132 87 147
rect 41 60 87 86
rect 521 198 567 209
rect 681 255 727 274
rect 361 60 407 83
rect 841 255 887 314
rect 841 198 887 209
rect 1001 255 1047 268
rect 681 60 727 81
rect 1161 255 1207 314
rect 1161 198 1207 209
rect 1321 255 1367 268
rect 1001 60 1047 81
rect 1481 255 1527 314
rect 1481 198 1527 209
rect 1641 254 1687 265
rect 1321 60 1367 81
rect 1801 255 1847 314
rect 1801 198 1847 209
rect 1641 60 1687 81
rect 0 -60 2016 60
<< labels >>
flabel metal1 s 0 724 2016 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2016 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 41 322 154 412 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 841 314 1847 396 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2016 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 2102 354
string MASKHINTS_PPLUS -86 354 2102 870
<< end >>
