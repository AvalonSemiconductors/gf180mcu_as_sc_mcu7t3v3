magic
tech gf180mcuD
magscale 1 5
timestamp 1751532423
<< nwell >>
rect -43 177 99 435
<< pwell >>
rect -43 -43 99 177
<< metal1 >>
rect 0 362 56 422
rect 0 -30 56 30
<< labels >>
flabel metal1 s 0 362 56 422 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -30 56 30 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 5 367 55 417 0 FreeSans 200 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 5 -25 55 25 0 FreeSans 200 0 0 0 VPW
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 56 392
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -8 -23 64 177
string MASKHINTS_PPLUS -8 177 64 415
<< end >>
