magic
tech gf180mcuD
magscale 1 10
timestamp 1764169223
<< nwell >>
rect -86 354 1766 870
<< pwell >>
rect -86 -86 1766 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 940 68 996 268
rect 1100 68 1156 268
rect 1260 68 1316 268
rect 1420 68 1476 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 940 440 996 716
rect 1100 440 1156 716
rect 1260 440 1316 716
rect 1420 440 1476 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 231 276 268
rect 172 185 201 231
rect 247 185 276 231
rect 172 68 276 185
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 231 596 268
rect 492 185 521 231
rect 567 185 596 231
rect 492 68 596 185
rect 652 127 740 268
rect 652 81 681 127
rect 727 81 740 127
rect 652 68 740 81
rect 796 255 940 268
rect 796 209 865 255
rect 911 209 940 255
rect 796 68 940 209
rect 996 152 1100 268
rect 996 106 1025 152
rect 1071 106 1100 152
rect 996 68 1100 106
rect 1156 233 1260 268
rect 1156 117 1185 233
rect 1231 117 1260 233
rect 1156 68 1260 117
rect 1316 255 1420 268
rect 1316 209 1345 255
rect 1391 209 1420 255
rect 1316 68 1420 209
rect 1476 152 1564 268
rect 1476 106 1505 152
rect 1551 106 1564 152
rect 1476 68 1564 106
<< pdiff >>
rect 28 624 116 716
rect 28 578 41 624
rect 87 578 116 624
rect 28 440 116 578
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 645 436 716
rect 332 599 361 645
rect 407 599 436 645
rect 332 440 436 599
rect 492 586 596 716
rect 492 540 521 586
rect 567 540 596 586
rect 492 440 596 540
rect 652 678 740 716
rect 652 632 681 678
rect 727 632 740 678
rect 652 440 740 632
rect 796 703 940 716
rect 796 657 865 703
rect 911 657 940 703
rect 796 440 940 657
rect 996 586 1100 716
rect 996 540 1025 586
rect 1071 540 1100 586
rect 996 440 1100 540
rect 1156 703 1260 716
rect 1156 657 1185 703
rect 1231 657 1260 703
rect 1156 440 1260 657
rect 1316 586 1420 716
rect 1316 453 1345 586
rect 1391 453 1420 586
rect 1316 440 1420 453
rect 1476 703 1564 716
rect 1476 657 1505 703
rect 1551 657 1564 703
rect 1476 440 1564 657
<< ndiffc >>
rect 41 81 87 127
rect 201 185 247 231
rect 361 81 407 127
rect 521 185 567 231
rect 681 81 727 127
rect 865 209 911 255
rect 1025 106 1071 152
rect 1185 117 1231 233
rect 1345 209 1391 255
rect 1505 106 1551 152
<< pdiffc >>
rect 41 578 87 624
rect 201 657 247 703
rect 361 599 407 645
rect 521 540 567 586
rect 681 632 727 678
rect 865 657 911 703
rect 1025 540 1071 586
rect 1185 657 1231 703
rect 1345 453 1391 586
rect 1505 657 1551 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 940 716 996 760
rect 1100 716 1156 760
rect 1260 716 1316 760
rect 1420 716 1476 760
rect 116 397 172 440
rect 276 397 332 440
rect 116 376 332 397
rect 116 330 129 376
rect 317 330 332 376
rect 116 316 332 330
rect 116 268 172 316
rect 276 268 332 316
rect 436 394 492 440
rect 596 394 652 440
rect 436 374 652 394
rect 436 328 452 374
rect 639 328 652 374
rect 436 313 652 328
rect 436 268 492 313
rect 596 268 652 313
rect 940 397 996 440
rect 1100 397 1156 440
rect 940 378 1156 397
rect 940 332 953 378
rect 1143 332 1156 378
rect 940 317 1156 332
rect 940 268 996 317
rect 1100 268 1156 317
rect 1260 393 1316 440
rect 1420 393 1476 440
rect 1260 377 1563 393
rect 1260 331 1503 377
rect 1549 331 1563 377
rect 1260 313 1563 331
rect 1260 268 1316 313
rect 1420 268 1476 313
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 940 24 996 68
rect 1100 24 1156 68
rect 1260 24 1316 68
rect 1420 24 1476 68
<< polycontact >>
rect 129 330 317 376
rect 452 328 639 374
rect 953 332 1143 378
rect 1503 331 1549 377
<< metal1 >>
rect 0 724 1680 844
rect 201 703 247 724
rect 865 703 911 724
rect 201 646 247 657
rect 41 624 87 646
rect 361 645 681 678
rect 87 599 361 600
rect 407 632 681 645
rect 727 632 738 678
rect 865 646 911 657
rect 1185 703 1231 724
rect 1185 646 1231 657
rect 1505 703 1551 724
rect 1505 646 1551 657
rect 87 578 407 599
rect 41 554 407 578
rect 505 540 521 586
rect 567 540 1025 586
rect 1071 540 1345 586
rect 930 397 998 494
rect 1391 453 1410 586
rect 124 376 317 397
rect 124 330 129 376
rect 124 316 317 330
rect 447 374 640 394
rect 447 328 452 374
rect 639 328 640 374
rect 447 313 640 328
rect 930 378 1156 397
rect 930 332 953 378
rect 1143 332 1156 378
rect 930 317 1156 332
rect 865 255 911 266
rect 186 185 201 231
rect 247 185 521 231
rect 567 185 819 231
rect 1345 255 1410 453
rect 1482 377 1628 393
rect 1482 331 1503 377
rect 1549 331 1628 377
rect 1482 313 1628 331
rect 911 233 1231 244
rect 911 209 1185 233
rect 865 198 1185 209
rect 773 152 819 185
rect 41 127 87 138
rect 41 60 87 81
rect 361 127 407 138
rect 361 60 407 81
rect 681 127 727 138
rect 773 106 1025 152
rect 1071 106 1083 152
rect 1391 209 1410 255
rect 1345 198 1410 209
rect 1231 117 1505 152
rect 1185 106 1505 117
rect 1551 106 1568 152
rect 681 60 727 81
rect 0 -60 1680 60
<< labels >>
flabel metal1 s 0 724 1680 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1680 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 124 316 317 397 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 447 313 640 394 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 930 317 1156 397 0 FreeSans 200 0 0 0 C
port 7 new signal input
flabel metal1 1345 198 1410 586 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel metal1 1482 313 1628 393 0 FreeSans 200 0 0 0 D
port 9 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1680 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1696 354
string MASKHINTS_PPLUS -16 354 1696 830
<< end >>
