magic
tech gf180mcuD
magscale 1 10
timestamp 1753172561
<< nwell >>
rect -86 354 1654 870
<< pwell >>
rect -86 -86 1654 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 884 68 940 268
rect 1044 68 1100 268
rect 1204 68 1260 268
rect 1364 68 1420 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 884 440 940 716
rect 1044 440 1100 716
rect 1204 440 1260 716
rect 1364 440 1420 716
<< ndiff >>
rect 28 230 116 268
rect 28 184 41 230
rect 87 184 116 230
rect 28 68 116 184
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 198 436 268
rect 332 152 361 198
rect 407 152 436 198
rect 332 68 436 152
rect 492 244 596 268
rect 492 198 521 244
rect 567 198 596 244
rect 492 68 596 198
rect 652 152 740 268
rect 652 106 681 152
rect 727 106 740 152
rect 652 68 740 106
rect 796 152 884 268
rect 796 106 809 152
rect 855 106 884 152
rect 796 68 884 106
rect 940 244 1044 268
rect 940 198 969 244
rect 1015 198 1044 244
rect 940 68 1044 198
rect 1100 152 1204 268
rect 1100 106 1129 152
rect 1175 106 1204 152
rect 1100 68 1204 106
rect 1260 255 1364 268
rect 1260 209 1289 255
rect 1335 209 1364 255
rect 1260 68 1364 209
rect 1420 152 1512 268
rect 1420 106 1449 152
rect 1495 106 1512 152
rect 1420 68 1512 106
<< pdiff >>
rect 28 703 116 716
rect 28 471 41 703
rect 87 471 116 703
rect 28 440 116 471
rect 172 667 276 716
rect 172 481 201 667
rect 247 481 276 667
rect 172 440 276 481
rect 332 703 436 716
rect 332 657 361 703
rect 407 657 436 703
rect 332 440 436 657
rect 492 667 596 716
rect 492 481 521 667
rect 567 481 596 667
rect 492 440 596 481
rect 652 703 884 716
rect 652 657 681 703
rect 855 657 884 703
rect 652 440 884 657
rect 940 598 1044 716
rect 940 552 969 598
rect 1015 552 1044 598
rect 940 440 1044 552
rect 1100 703 1204 716
rect 1100 657 1129 703
rect 1175 657 1204 703
rect 1100 440 1204 657
rect 1260 592 1364 716
rect 1260 546 1289 592
rect 1335 546 1364 592
rect 1260 440 1364 546
rect 1420 703 1512 716
rect 1420 453 1449 703
rect 1495 453 1512 703
rect 1420 440 1512 453
<< ndiffc >>
rect 41 184 87 230
rect 201 81 247 127
rect 361 152 407 198
rect 521 198 567 244
rect 681 106 727 152
rect 809 106 855 152
rect 969 198 1015 244
rect 1129 106 1175 152
rect 1289 209 1335 255
rect 1449 106 1495 152
<< pdiffc >>
rect 41 471 87 703
rect 201 481 247 667
rect 361 657 407 703
rect 521 481 567 667
rect 681 657 855 703
rect 969 552 1015 598
rect 1129 657 1175 703
rect 1289 546 1335 592
rect 1449 453 1495 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 884 716 940 760
rect 1044 716 1100 760
rect 1204 716 1260 760
rect 1364 716 1420 760
rect 116 394 172 440
rect 276 394 332 440
rect 75 380 332 394
rect 436 391 492 440
rect 596 391 652 440
rect 884 394 940 440
rect 75 334 88 380
rect 285 334 332 380
rect 75 317 332 334
rect 116 268 172 317
rect 276 268 332 317
rect 395 375 652 391
rect 395 329 408 375
rect 639 329 652 375
rect 395 314 652 329
rect 836 378 940 394
rect 1044 378 1100 440
rect 1204 394 1260 440
rect 836 332 850 378
rect 896 332 1100 378
rect 836 317 940 332
rect 436 268 492 314
rect 596 268 652 314
rect 884 268 940 317
rect 1044 268 1100 332
rect 1156 382 1260 394
rect 1364 382 1420 440
rect 1156 378 1420 382
rect 1156 332 1174 378
rect 1220 332 1420 378
rect 1156 328 1420 332
rect 1156 317 1260 328
rect 1204 268 1260 317
rect 1364 268 1420 328
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 884 24 940 68
rect 1044 24 1100 68
rect 1204 24 1260 68
rect 1364 24 1420 68
<< polycontact >>
rect 88 334 285 380
rect 408 329 639 375
rect 850 332 896 378
rect 1174 332 1220 378
<< metal1 >>
rect 0 724 1568 844
rect 41 703 87 724
rect 361 703 407 724
rect 41 460 87 471
rect 201 667 247 678
rect 681 703 855 724
rect 361 646 407 657
rect 521 667 567 678
rect 247 481 521 516
rect 681 646 855 657
rect 1129 703 1175 724
rect 1129 646 1175 657
rect 1449 703 1495 724
rect 969 598 1015 609
rect 567 552 969 575
rect 1289 592 1335 609
rect 1015 552 1289 575
rect 567 546 1289 552
rect 567 529 1335 546
rect 1289 512 1335 529
rect 201 470 567 481
rect 75 380 285 394
rect 75 334 88 380
rect 75 317 285 334
rect 395 375 652 391
rect 395 329 408 375
rect 639 329 652 375
rect 395 314 652 329
rect 836 378 916 483
rect 836 332 850 378
rect 896 332 916 378
rect 836 317 916 332
rect 1156 378 1236 483
rect 1156 332 1174 378
rect 1220 332 1236 378
rect 1156 317 1236 332
rect 1289 255 1375 512
rect 1449 430 1495 453
rect 41 230 87 241
rect 87 198 407 230
rect 471 198 521 244
rect 567 198 969 244
rect 1015 198 1026 244
rect 1335 209 1375 255
rect 1289 198 1375 209
rect 87 184 361 198
rect 41 173 87 184
rect 201 127 247 138
rect 361 106 681 152
rect 727 106 738 152
rect 798 106 809 152
rect 855 106 1129 152
rect 1175 106 1449 152
rect 1495 106 1506 152
rect 201 60 247 81
rect 0 -60 1568 60
<< labels >>
flabel metal1 s 0 724 1568 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1568 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 75 317 285 394 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 395 314 652 391 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 836 317 916 483 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 1156 317 1236 483 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel metal1 1289 198 1375 512 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1584 354
string MASKHINTS_PPLUS -16 354 1584 830
<< end >>
