magic
tech gf180mcuD
magscale 1 10
timestamp 1753277880
<< nwell >>
rect -86 354 1990 870
<< pwell >>
rect -86 -86 1990 354
<< nmos >>
rect 116 68 172 268
rect 388 68 444 268
rect 500 68 556 268
rect 804 68 860 268
rect 984 68 1040 268
rect 1144 68 1200 268
rect 1314 68 1370 268
rect 1474 68 1530 268
rect 1634 68 1690 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 500 440 556 716
rect 700 440 756 716
rect 984 440 1040 716
rect 1144 440 1200 716
rect 1314 440 1370 716
rect 1474 440 1530 716
rect 1634 440 1690 716
<< ndiff >>
rect 28 255 116 268
rect 28 209 41 255
rect 87 209 116 255
rect 28 68 116 209
rect 172 127 388 268
rect 172 81 201 127
rect 247 81 388 127
rect 172 68 388 81
rect 444 68 500 268
rect 556 255 804 268
rect 556 209 585 255
rect 631 209 804 255
rect 556 68 804 209
rect 860 255 984 268
rect 860 209 909 255
rect 955 209 984 255
rect 860 68 984 209
rect 1040 127 1144 268
rect 1040 81 1069 127
rect 1115 81 1144 127
rect 1040 68 1144 81
rect 1200 255 1314 268
rect 1200 209 1239 255
rect 1285 209 1314 255
rect 1200 68 1314 209
rect 1370 255 1474 268
rect 1370 81 1399 255
rect 1445 81 1474 255
rect 1370 68 1474 81
rect 1530 255 1634 268
rect 1530 209 1559 255
rect 1605 209 1634 255
rect 1530 68 1634 209
rect 1690 255 1802 268
rect 1690 81 1719 255
rect 1765 81 1802 255
rect 1690 68 1802 81
<< pdiff >>
rect 28 667 116 716
rect 28 453 41 667
rect 87 453 116 667
rect 28 440 116 453
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 440 500 716
rect 556 599 700 716
rect 556 553 585 599
rect 631 553 700 599
rect 556 440 700 553
rect 756 507 984 716
rect 756 461 785 507
rect 831 461 984 507
rect 756 440 984 461
rect 1040 703 1144 716
rect 1040 657 1069 703
rect 1115 657 1144 703
rect 1040 440 1144 657
rect 1200 667 1314 716
rect 1200 453 1239 667
rect 1285 453 1314 667
rect 1200 440 1314 453
rect 1370 703 1474 716
rect 1370 453 1399 703
rect 1445 453 1474 703
rect 1370 440 1474 453
rect 1530 667 1634 716
rect 1530 453 1559 667
rect 1605 453 1634 667
rect 1530 440 1634 453
rect 1690 703 1796 716
rect 1690 453 1719 703
rect 1765 453 1796 703
rect 1690 440 1796 453
<< ndiffc >>
rect 41 209 87 255
rect 201 81 247 127
rect 585 209 631 255
rect 909 209 955 255
rect 1069 81 1115 127
rect 1239 209 1285 255
rect 1399 81 1445 255
rect 1559 209 1605 255
rect 1719 81 1765 255
<< pdiffc >>
rect 41 453 87 667
rect 201 657 247 703
rect 585 553 631 599
rect 785 461 831 507
rect 1069 657 1115 703
rect 1239 453 1285 667
rect 1399 453 1445 703
rect 1559 453 1605 667
rect 1719 453 1765 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 500 716 556 760
rect 700 716 756 760
rect 984 716 1040 760
rect 1144 716 1200 760
rect 1314 716 1370 760
rect 1474 716 1530 760
rect 1634 716 1690 760
rect 116 420 172 440
rect 276 420 332 440
rect 116 375 332 420
rect 500 388 556 440
rect 700 388 756 440
rect 984 392 1040 440
rect 1144 392 1200 440
rect 1314 392 1370 440
rect 116 329 133 375
rect 179 374 332 375
rect 380 375 452 388
rect 179 329 192 374
rect 116 316 192 329
rect 380 329 393 375
rect 439 329 452 375
rect 380 316 452 329
rect 500 375 636 388
rect 500 329 577 375
rect 623 329 636 375
rect 500 316 636 329
rect 684 375 756 388
rect 684 329 697 375
rect 743 329 756 375
rect 684 316 756 329
rect 804 375 876 388
rect 804 329 817 375
rect 863 329 876 375
rect 804 316 876 329
rect 984 379 1060 392
rect 984 333 1001 379
rect 1047 333 1060 379
rect 984 320 1060 333
rect 1134 379 1370 392
rect 1474 383 1530 440
rect 1634 383 1690 440
rect 1474 379 1690 383
rect 1134 333 1147 379
rect 1193 333 1690 379
rect 1134 332 1690 333
rect 1134 320 1370 332
rect 116 268 172 316
rect 388 268 444 316
rect 500 268 556 316
rect 804 268 860 316
rect 984 268 1040 320
rect 1144 268 1200 320
rect 1314 268 1370 320
rect 1474 268 1530 332
rect 1634 268 1690 332
rect 116 24 172 68
rect 388 24 444 68
rect 500 24 556 68
rect 804 24 860 68
rect 984 24 1040 68
rect 1144 24 1200 68
rect 1314 24 1370 68
rect 1474 24 1530 68
rect 1634 24 1690 68
<< polycontact >>
rect 133 329 179 375
rect 393 329 439 375
rect 577 329 623 375
rect 697 329 743 375
rect 817 329 863 375
rect 1001 333 1047 379
rect 1147 333 1193 379
<< metal1 >>
rect 0 724 1904 844
rect 201 703 247 724
rect 41 667 87 678
rect 201 646 247 657
rect 1069 703 1115 724
rect 1399 703 1445 724
rect 1069 646 1115 657
rect 1239 667 1310 678
rect 139 577 151 629
rect 485 553 585 599
rect 631 553 1193 599
rect 387 537 439 549
rect 41 268 87 453
rect 133 485 387 531
rect 133 375 208 485
rect 387 473 439 485
rect 179 329 208 375
rect 133 318 208 329
rect 393 375 439 400
rect 393 268 439 329
rect 41 255 439 268
rect 87 222 439 255
rect 485 255 531 553
rect 577 461 785 507
rect 831 461 955 507
rect 577 375 623 461
rect 577 313 623 329
rect 684 403 743 415
rect 684 351 688 403
rect 740 375 743 403
rect 684 329 697 351
rect 684 316 743 329
rect 817 375 863 388
rect 485 209 585 255
rect 631 209 642 255
rect 688 247 740 249
rect 817 247 863 329
rect 688 237 863 247
rect 41 198 87 209
rect 740 201 863 237
rect 909 255 955 461
rect 1001 379 1088 402
rect 1147 392 1193 553
rect 1047 333 1088 379
rect 1001 320 1088 333
rect 1134 379 1193 392
rect 1134 333 1147 379
rect 1134 320 1193 333
rect 1285 453 1310 667
rect 1239 379 1310 453
rect 1719 703 1765 724
rect 1399 435 1445 453
rect 1559 667 1619 678
rect 1605 453 1619 667
rect 1559 379 1619 453
rect 1719 434 1765 453
rect 1239 333 1619 379
rect 909 196 955 209
rect 1239 255 1310 333
rect 1285 209 1310 255
rect 1239 198 1310 209
rect 1399 255 1445 275
rect 688 173 740 185
rect 201 127 247 138
rect 201 60 247 81
rect 1069 127 1115 138
rect 1069 60 1115 81
rect 1559 255 1619 333
rect 1605 209 1619 255
rect 1559 198 1619 209
rect 1719 255 1765 275
rect 1399 60 1445 81
rect 1719 60 1765 81
rect 0 -60 1904 60
<< via1 >>
rect 87 577 139 629
rect 387 485 439 537
rect 688 375 740 403
rect 688 351 697 375
rect 697 351 740 375
rect 688 185 740 237
<< metal2 >>
rect 75 631 142 632
rect 263 631 742 651
rect 75 629 742 631
rect 75 577 87 629
rect 139 595 742 629
rect 139 577 319 595
rect 75 575 319 577
rect 75 574 142 575
rect 375 537 451 539
rect 375 485 387 537
rect 439 485 451 537
rect 375 473 451 485
rect 393 238 449 473
rect 686 406 742 595
rect 684 403 743 406
rect 684 351 688 403
rect 740 351 743 403
rect 684 339 743 351
rect 682 238 746 249
rect 393 237 746 238
rect 393 185 688 237
rect 740 185 746 237
rect 393 182 746 185
rect 682 173 746 182
<< labels >>
flabel metal1 s 0 724 1904 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1904 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 1001 320 1088 402 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel metal1 133 318 208 531 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 1239 198 1310 678 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel metal1 1559 198 1619 678 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1904 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1920 354
string MASKHINTS_PPLUS -16 354 1920 830
<< end >>
