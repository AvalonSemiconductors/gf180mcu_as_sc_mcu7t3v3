magic
tech gf180mcuD
magscale 1 10
timestamp 1764156381
<< nwell >>
rect -86 354 2886 870
<< pwell >>
rect -86 -86 2886 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
rect 1396 68 1452 268
rect 1556 68 1612 268
rect 1716 68 1772 268
rect 1876 68 1932 268
rect 2036 68 2092 268
rect 2196 68 2252 268
rect 2356 68 2412 268
rect 2516 68 2572 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1396 440 1452 716
rect 1556 440 1612 716
rect 1716 440 1772 716
rect 1876 440 1932 716
rect 2036 440 2092 716
rect 2196 440 2252 716
rect 2356 440 2412 716
rect 2516 440 2572 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 218 276 268
rect 172 172 201 218
rect 247 172 276 218
rect 172 68 276 172
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 163 596 268
rect 492 117 521 163
rect 567 117 596 163
rect 492 68 596 117
rect 652 244 756 268
rect 652 198 681 244
rect 727 198 756 244
rect 652 68 756 198
rect 812 152 916 268
rect 812 106 841 152
rect 887 106 916 152
rect 812 68 916 106
rect 972 244 1076 268
rect 972 198 1001 244
rect 1047 198 1076 244
rect 972 68 1076 198
rect 1132 152 1236 268
rect 1132 106 1161 152
rect 1207 106 1236 152
rect 1132 68 1236 106
rect 1292 127 1396 268
rect 1292 81 1321 127
rect 1367 81 1396 127
rect 1292 68 1396 81
rect 1452 244 1556 268
rect 1452 198 1481 244
rect 1527 198 1556 244
rect 1452 68 1556 198
rect 1612 127 1716 268
rect 1612 81 1641 127
rect 1687 81 1716 127
rect 1612 68 1716 81
rect 1772 244 1876 268
rect 1772 198 1801 244
rect 1847 198 1876 244
rect 1772 68 1876 198
rect 1932 127 2036 268
rect 1932 81 1961 127
rect 2007 81 2036 127
rect 1932 68 2036 81
rect 2092 244 2196 268
rect 2092 198 2121 244
rect 2167 198 2196 244
rect 2092 68 2196 198
rect 2252 127 2356 268
rect 2252 81 2281 127
rect 2327 81 2356 127
rect 2252 68 2356 81
rect 2412 244 2516 268
rect 2412 198 2441 244
rect 2487 198 2516 244
rect 2412 68 2516 198
rect 2572 127 2660 268
rect 2572 81 2601 127
rect 2647 81 2660 127
rect 2572 68 2660 81
<< pdiff >>
rect 28 644 116 716
rect 28 598 41 644
rect 87 598 116 644
rect 28 440 116 598
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 600 436 716
rect 332 554 361 600
rect 407 554 436 600
rect 332 440 436 554
rect 492 703 596 716
rect 492 657 521 703
rect 567 657 596 703
rect 492 440 596 657
rect 652 600 756 716
rect 652 554 681 600
rect 727 554 756 600
rect 652 440 756 554
rect 812 703 916 716
rect 812 657 841 703
rect 887 657 916 703
rect 812 440 916 657
rect 972 600 1076 716
rect 972 554 1001 600
rect 1047 554 1076 600
rect 972 440 1076 554
rect 1132 703 1236 716
rect 1132 657 1161 703
rect 1207 657 1236 703
rect 1132 440 1236 657
rect 1292 611 1396 716
rect 1292 565 1321 611
rect 1367 565 1396 611
rect 1292 440 1396 565
rect 1452 499 1556 716
rect 1452 453 1481 499
rect 1527 453 1556 499
rect 1452 440 1556 453
rect 1612 678 1716 716
rect 1612 632 1641 678
rect 1687 632 1716 678
rect 1612 440 1716 632
rect 1772 440 1876 716
rect 1932 595 2036 716
rect 1932 549 1961 595
rect 2007 549 2036 595
rect 1932 440 2036 549
rect 2092 499 2196 716
rect 2092 453 2121 499
rect 2167 453 2196 499
rect 2092 440 2196 453
rect 2252 595 2356 716
rect 2252 549 2281 595
rect 2327 549 2356 595
rect 2252 440 2356 549
rect 2412 440 2516 716
rect 2572 654 2660 716
rect 2572 608 2601 654
rect 2647 608 2660 654
rect 2572 440 2660 608
<< ndiffc >>
rect 41 81 87 127
rect 201 172 247 218
rect 361 81 407 127
rect 521 117 567 163
rect 681 198 727 244
rect 841 106 887 152
rect 1001 198 1047 244
rect 1161 106 1207 152
rect 1321 81 1367 127
rect 1481 198 1527 244
rect 1641 81 1687 127
rect 1801 198 1847 244
rect 1961 81 2007 127
rect 2121 198 2167 244
rect 2281 81 2327 127
rect 2441 198 2487 244
rect 2601 81 2647 127
<< pdiffc >>
rect 41 598 87 644
rect 201 657 247 703
rect 361 554 407 600
rect 521 657 567 703
rect 681 554 727 600
rect 841 657 887 703
rect 1001 554 1047 600
rect 1161 657 1207 703
rect 1321 565 1367 611
rect 1481 453 1527 499
rect 1641 632 1687 678
rect 1961 549 2007 595
rect 2121 453 2167 499
rect 2281 549 2327 595
rect 2601 608 2647 654
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1396 716 1452 760
rect 1556 716 1612 760
rect 1716 716 1772 760
rect 1876 716 1932 760
rect 2036 716 2092 760
rect 2196 716 2252 760
rect 2356 716 2412 760
rect 2516 716 2572 760
rect 116 393 172 440
rect 276 393 332 440
rect 436 393 492 440
rect 116 373 492 393
rect 116 327 129 373
rect 479 327 492 373
rect 116 314 492 327
rect 116 268 172 314
rect 276 268 332 314
rect 436 268 492 314
rect 596 392 652 440
rect 756 392 812 440
rect 916 392 972 440
rect 1076 392 1132 440
rect 596 374 1132 392
rect 1236 388 1292 440
rect 1396 391 1452 440
rect 1556 391 1612 440
rect 1716 391 1772 440
rect 596 327 609 374
rect 1113 327 1132 374
rect 596 304 1132 327
rect 1228 376 1300 388
rect 1228 330 1241 376
rect 1287 330 1300 376
rect 1228 318 1300 330
rect 1396 374 1772 391
rect 1396 327 1409 374
rect 1759 327 1772 374
rect 596 268 652 304
rect 756 268 812 304
rect 916 268 972 304
rect 1076 268 1132 304
rect 1236 268 1292 318
rect 1396 313 1772 327
rect 1396 268 1452 313
rect 1556 268 1612 313
rect 1716 268 1772 313
rect 1876 392 1932 440
rect 2036 392 2092 440
rect 2196 392 2252 440
rect 2356 392 2412 440
rect 1876 379 2412 392
rect 2516 388 2572 440
rect 1876 333 1889 379
rect 2396 333 2412 379
rect 1876 320 2412 333
rect 1876 268 1932 320
rect 2036 268 2092 320
rect 2196 268 2252 320
rect 2356 268 2412 320
rect 2508 376 2580 388
rect 2508 330 2521 376
rect 2567 330 2580 376
rect 2508 318 2580 330
rect 2516 268 2572 318
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1396 24 1452 68
rect 1556 24 1612 68
rect 1716 24 1772 68
rect 1876 24 1932 68
rect 2036 24 2092 68
rect 2196 24 2252 68
rect 2356 24 2412 68
rect 2516 24 2572 68
<< polycontact >>
rect 129 327 479 373
rect 609 327 1113 374
rect 1241 330 1287 376
rect 1409 327 1759 374
rect 1889 333 2396 379
rect 2521 330 2567 376
<< metal1 >>
rect 0 724 2800 844
rect 201 703 247 724
rect 41 644 87 678
rect 201 646 247 657
rect 521 703 567 724
rect 521 646 567 657
rect 841 703 887 724
rect 841 646 887 657
rect 1161 703 1207 724
rect 1161 646 1207 657
rect 1321 632 1641 678
rect 1687 657 1719 678
rect 1321 611 1367 632
rect 87 598 361 600
rect 41 554 361 598
rect 407 554 681 600
rect 727 554 1001 600
rect 1047 565 1321 600
rect 1641 605 1656 632
rect 1708 605 1719 657
rect 1641 591 1719 605
rect 2583 654 2647 678
rect 2583 650 2601 654
rect 2583 598 2588 650
rect 2640 598 2647 608
rect 1047 554 1367 565
rect 1950 549 1961 595
rect 2007 549 2281 595
rect 2327 549 2474 595
rect 2583 586 2647 598
rect 2428 540 2474 549
rect 425 443 1287 489
rect 1470 453 1481 499
rect 1527 494 1538 499
rect 2110 494 2121 499
rect 1527 453 2121 494
rect 2167 453 2178 499
rect 2428 494 2695 540
rect 1470 448 2178 453
rect 425 395 492 443
rect 116 373 492 395
rect 116 327 129 373
rect 479 327 492 373
rect 116 315 492 327
rect 596 374 1113 392
rect 596 327 609 374
rect 596 313 1113 327
rect 1241 376 1287 443
rect 1241 314 1287 330
rect 1396 374 1777 391
rect 1396 327 1409 374
rect 1759 369 1777 374
rect 1396 317 1713 327
rect 1765 317 1777 369
rect 1876 379 2403 388
rect 1876 333 1889 379
rect 2396 333 2403 379
rect 1876 320 2403 333
rect 2497 378 2580 388
rect 2497 326 2518 378
rect 2570 326 2580 378
rect 2497 318 2580 326
rect 1396 313 1777 317
rect 2626 244 2695 494
rect 201 218 567 230
rect 247 184 567 218
rect 670 198 681 244
rect 727 198 1001 244
rect 1047 198 1481 244
rect 1527 198 1801 244
rect 1847 198 2121 244
rect 2167 198 2441 244
rect 2487 198 2695 244
rect 201 158 247 172
rect 521 163 567 184
rect 41 127 87 138
rect 41 60 87 81
rect 361 127 407 138
rect 567 117 841 152
rect 521 106 841 117
rect 887 106 1161 152
rect 1207 106 1219 152
rect 1321 127 1367 138
rect 361 60 407 81
rect 1321 60 1367 81
rect 1641 127 1687 138
rect 1641 60 1687 81
rect 1961 127 2007 138
rect 1961 60 2007 81
rect 2281 127 2327 138
rect 2281 60 2327 81
rect 2601 127 2647 138
rect 2601 60 2647 81
rect 0 -60 2800 60
<< via1 >>
rect 1656 632 1687 657
rect 1687 632 1708 657
rect 1656 605 1708 632
rect 2588 608 2601 650
rect 2601 608 2640 650
rect 2588 598 2640 608
rect 1713 327 1759 369
rect 1759 327 1765 369
rect 1713 317 1765 327
rect 2518 376 2570 378
rect 2518 330 2521 376
rect 2521 330 2567 376
rect 2567 330 2570 376
rect 2518 326 2570 330
<< metal2 >>
rect 1644 657 1720 661
rect 1644 605 1656 657
rect 1708 647 1720 657
rect 2576 650 2645 662
rect 2576 647 2588 650
rect 1708 605 2588 647
rect 1644 598 2588 605
rect 2640 598 2645 650
rect 1644 591 2645 598
rect 2576 586 2645 591
rect 1711 369 1777 381
rect 1711 317 1713 369
rect 1765 317 1777 369
rect 1711 264 1777 317
rect 2516 378 2572 390
rect 2516 326 2518 378
rect 2570 326 2572 378
rect 2516 264 2572 326
rect 1711 208 2572 264
<< labels >>
flabel metal1 s 0 724 2800 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2800 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 116 315 492 395 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 596 313 1113 392 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 1396 313 1713 391 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 1876 320 2403 388 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel metal1 2626 198 2695 540 0 FreeSans 200 0 0 0 Y
port 9 new signal output
<< properties >>
string FIXED_BBOX 0 0 2800 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 2816 354
string MASKHINTS_PPLUS -16 354 2816 830
<< end >>
