magic
tech gf180mcuD
magscale 1 10
timestamp 1758891449
<< nwell >>
rect -86 354 3110 870
<< pwell >>
rect -86 -86 3110 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 573 68 629 268
rect 797 68 853 268
rect 1203 68 1259 268
rect 1315 68 1371 268
rect 1475 68 1531 268
rect 1653 68 1709 268
rect 1959 68 2015 268
rect 2187 68 2243 268
rect 2347 68 2403 268
rect 2657 68 2713 268
rect 2817 68 2873 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 678 440 735 716
rect 797 440 853 716
rect 1007 440 1064 716
rect 1315 440 1371 716
rect 1475 440 1531 716
rect 1772 440 1828 716
rect 2072 440 2128 716
rect 2187 440 2243 716
rect 2347 440 2403 716
rect 2657 440 2713 716
rect 2817 440 2873 716
<< ndiff >>
rect 28 255 116 268
rect 28 209 41 255
rect 87 209 116 255
rect 28 68 116 209
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 255 429 268
rect 332 209 361 255
rect 407 209 429 255
rect 332 68 429 209
rect 485 127 573 268
rect 485 81 498 127
rect 544 81 573 127
rect 485 68 573 81
rect 629 68 797 268
rect 853 255 1203 268
rect 853 209 932 255
rect 978 209 1203 255
rect 853 68 1203 209
rect 1259 68 1315 268
rect 1371 127 1475 268
rect 1371 81 1400 127
rect 1446 81 1475 127
rect 1371 68 1475 81
rect 1531 255 1653 268
rect 1531 209 1560 255
rect 1606 209 1653 255
rect 1531 68 1653 209
rect 1709 255 1959 268
rect 1709 209 1884 255
rect 1930 209 1959 255
rect 1709 68 1959 209
rect 2015 68 2187 268
rect 2243 127 2347 268
rect 2243 81 2272 127
rect 2318 81 2347 127
rect 2243 68 2347 81
rect 2403 255 2513 268
rect 2403 209 2454 255
rect 2500 209 2513 255
rect 2403 68 2513 209
rect 2569 255 2657 268
rect 2569 81 2582 255
rect 2628 81 2657 255
rect 2569 68 2657 81
rect 2713 255 2817 268
rect 2713 209 2742 255
rect 2788 209 2817 255
rect 2713 68 2817 209
rect 2873 255 2996 268
rect 2873 81 2902 255
rect 2948 81 2996 255
rect 2873 68 2996 81
<< pdiff >>
rect 28 587 116 716
rect 28 541 41 587
rect 87 541 116 587
rect 28 440 116 541
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 667 429 716
rect 332 501 361 667
rect 407 501 429 667
rect 332 440 429 501
rect 485 703 678 716
rect 485 657 498 703
rect 544 657 678 703
rect 485 440 678 657
rect 735 440 797 716
rect 853 499 1007 716
rect 853 453 932 499
rect 978 453 1007 499
rect 853 440 1007 453
rect 1064 440 1315 716
rect 1371 703 1475 716
rect 1371 657 1400 703
rect 1446 657 1475 703
rect 1371 440 1475 657
rect 1531 499 1772 716
rect 1531 453 1560 499
rect 1606 453 1772 499
rect 1531 440 1772 453
rect 1828 499 2072 716
rect 1828 453 1884 499
rect 1930 453 2072 499
rect 1828 440 2072 453
rect 2128 440 2187 716
rect 2243 703 2347 716
rect 2243 657 2272 703
rect 2318 657 2347 703
rect 2243 440 2347 657
rect 2403 667 2513 716
rect 2403 453 2454 667
rect 2500 453 2513 667
rect 2403 440 2513 453
rect 2569 703 2657 716
rect 2569 453 2582 703
rect 2628 453 2657 703
rect 2569 440 2657 453
rect 2713 499 2817 716
rect 2713 453 2742 499
rect 2788 453 2817 499
rect 2713 440 2817 453
rect 2873 703 2996 716
rect 2873 453 2902 703
rect 2948 453 2996 703
rect 2873 440 2996 453
<< ndiffc >>
rect 41 209 87 255
rect 201 81 247 127
rect 361 209 407 255
rect 498 81 544 127
rect 932 209 978 255
rect 1400 81 1446 127
rect 1560 209 1606 255
rect 1884 209 1930 255
rect 2272 81 2318 127
rect 2454 209 2500 255
rect 2582 81 2628 255
rect 2742 209 2788 255
rect 2902 81 2948 255
<< pdiffc >>
rect 41 541 87 587
rect 201 657 247 703
rect 361 501 407 667
rect 498 657 544 703
rect 932 453 978 499
rect 1400 657 1446 703
rect 1560 453 1606 499
rect 1884 453 1930 499
rect 2272 657 2318 703
rect 2454 453 2500 667
rect 2582 453 2628 703
rect 2742 453 2788 499
rect 2902 453 2948 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 678 716 735 760
rect 797 716 853 760
rect 1007 716 1064 760
rect 1315 716 1371 760
rect 1475 716 1531 760
rect 1772 716 1828 760
rect 2072 716 2128 760
rect 2187 716 2243 760
rect 2347 716 2403 760
rect 2657 716 2713 760
rect 2817 716 2873 760
rect 116 394 172 440
rect 100 379 172 394
rect 276 420 332 440
rect 276 407 509 420
rect 276 393 450 407
rect 100 333 113 379
rect 159 333 172 379
rect 100 320 172 333
rect 116 268 172 320
rect 222 378 450 393
rect 222 332 235 378
rect 281 375 450 378
rect 281 332 332 375
rect 437 361 450 375
rect 496 361 509 407
rect 678 406 735 440
rect 437 348 509 361
rect 677 393 749 406
rect 222 319 332 332
rect 276 268 332 319
rect 557 347 629 360
rect 557 301 570 347
rect 616 301 629 347
rect 677 347 690 393
rect 736 347 749 393
rect 677 334 749 347
rect 797 398 853 440
rect 1007 398 1064 440
rect 1315 398 1371 440
rect 797 385 869 398
rect 797 339 810 385
rect 856 339 869 385
rect 557 288 629 301
rect 573 268 629 288
rect 797 326 869 339
rect 1007 385 1083 398
rect 1007 339 1024 385
rect 1070 339 1083 385
rect 1007 326 1083 339
rect 1195 385 1267 398
rect 1195 339 1208 385
rect 1254 339 1267 385
rect 1195 326 1267 339
rect 1315 385 1387 398
rect 1475 397 1531 440
rect 1772 397 1828 440
rect 2072 397 2128 440
rect 2187 397 2243 440
rect 1315 339 1328 385
rect 1374 339 1387 385
rect 1315 326 1387 339
rect 1446 384 1531 397
rect 1446 338 1460 384
rect 1506 338 1531 384
rect 797 268 853 326
rect 1203 268 1259 326
rect 1315 268 1371 326
rect 1446 325 1531 338
rect 1652 384 1724 397
rect 1652 338 1665 384
rect 1711 338 1724 384
rect 1652 325 1724 338
rect 1772 384 1844 397
rect 1772 338 1785 384
rect 1831 371 1844 384
rect 2063 384 2139 397
rect 1831 338 2015 371
rect 1772 325 2015 338
rect 2063 338 2078 384
rect 2124 338 2139 384
rect 2063 325 2139 338
rect 2187 384 2263 397
rect 2187 338 2202 384
rect 2248 338 2263 384
rect 2187 325 2263 338
rect 2347 396 2403 440
rect 2657 396 2713 440
rect 2817 396 2873 440
rect 2347 383 2423 396
rect 2347 337 2362 383
rect 2408 337 2423 383
rect 1475 268 1531 325
rect 1653 268 1709 325
rect 1959 268 2015 325
rect 2187 268 2243 325
rect 2347 324 2423 337
rect 2471 383 2873 396
rect 2471 337 2484 383
rect 2530 337 2873 383
rect 2471 324 2873 337
rect 2347 268 2403 324
rect 2657 268 2713 324
rect 2817 268 2873 324
rect 116 24 172 68
rect 276 24 332 68
rect 573 24 629 68
rect 797 24 853 68
rect 1203 24 1259 68
rect 1315 24 1371 68
rect 1475 24 1531 68
rect 1653 24 1709 68
rect 1959 24 2015 68
rect 2187 24 2243 68
rect 2347 24 2403 68
rect 2657 24 2713 68
rect 2817 24 2873 68
<< polycontact >>
rect 113 333 159 379
rect 235 332 281 378
rect 450 361 496 407
rect 570 301 616 347
rect 690 347 736 393
rect 810 339 856 385
rect 1024 339 1070 385
rect 1208 339 1254 385
rect 1328 339 1374 385
rect 1460 338 1506 384
rect 1665 338 1711 384
rect 1785 338 1831 384
rect 2078 338 2124 384
rect 2202 338 2248 384
rect 2362 337 2408 383
rect 2484 337 2530 383
<< metal1 >>
rect 0 724 3024 844
rect 201 703 247 724
rect 498 703 544 724
rect 201 646 247 657
rect 358 667 407 678
rect 41 587 89 599
rect 87 541 267 587
rect 41 530 89 541
rect 25 379 172 412
rect 25 333 113 379
rect 159 333 172 379
rect 25 320 172 333
rect 221 397 267 541
rect 358 501 361 667
rect 1400 703 1446 724
rect 498 646 544 657
rect 594 632 1241 678
rect 1400 646 1446 657
rect 2272 703 2318 724
rect 2582 703 2628 724
rect 594 600 640 632
rect 407 554 640 600
rect 358 490 407 501
rect 221 378 281 397
rect 221 332 235 378
rect 221 321 281 332
rect 41 255 87 266
rect 221 255 267 321
rect 358 310 404 490
rect 450 409 736 455
rect 450 407 496 409
rect 450 344 496 361
rect 690 393 736 409
rect 570 347 616 358
rect 358 256 407 310
rect 570 256 616 301
rect 87 209 267 255
rect 350 255 616 256
rect 350 209 361 255
rect 407 209 616 255
rect 41 198 87 209
rect 690 152 736 347
rect 797 385 886 586
rect 797 339 810 385
rect 856 339 886 385
rect 797 326 886 339
rect 932 499 978 510
rect 932 280 978 453
rect 1024 385 1070 632
rect 1185 618 1241 632
rect 1185 606 1261 618
rect 1185 554 1197 606
rect 1249 554 1261 606
rect 1185 551 1261 554
rect 1664 601 2124 647
rect 2272 646 2318 657
rect 2454 667 2500 678
rect 1024 326 1070 339
rect 1116 459 1506 505
rect 1116 280 1162 459
rect 1209 398 1265 405
rect 932 255 1162 280
rect 978 234 1162 255
rect 1208 393 1265 398
rect 1208 385 1209 393
rect 1261 341 1265 393
rect 1254 339 1265 341
rect 1208 329 1265 339
rect 1325 385 1377 398
rect 1325 339 1328 385
rect 1374 339 1377 385
rect 932 198 978 209
rect 1208 152 1254 329
rect 1325 328 1377 339
rect 1331 244 1377 328
rect 1460 384 1506 459
rect 1460 325 1506 338
rect 1560 499 1606 510
rect 1560 255 1606 453
rect 1664 397 1710 601
rect 1884 499 1930 510
rect 1652 393 1728 397
rect 1652 341 1664 393
rect 1716 341 1728 393
rect 1652 338 1665 341
rect 1711 338 1728 341
rect 1652 319 1728 338
rect 1774 392 1838 405
rect 1774 384 1786 392
rect 1774 338 1785 384
rect 1831 338 1838 340
rect 1774 312 1838 338
rect 1331 209 1560 244
rect 1331 198 1606 209
rect 1884 255 1930 453
rect 2078 384 2124 601
rect 2078 325 2124 338
rect 2202 454 2454 500
rect 2202 384 2248 454
rect 2454 396 2500 453
rect 2902 703 2948 724
rect 2582 429 2628 453
rect 2723 499 2809 510
rect 2723 453 2742 499
rect 2788 453 2809 499
rect 2202 325 2248 338
rect 2362 383 2408 396
rect 2362 230 2408 337
rect 1930 209 2408 230
rect 1884 184 2408 209
rect 2454 383 2530 396
rect 2454 337 2484 383
rect 2454 324 2530 337
rect 2454 255 2500 324
rect 2454 198 2500 209
rect 2582 255 2628 278
rect 201 127 247 138
rect 201 60 247 81
rect 498 127 544 138
rect 690 106 1254 152
rect 1400 127 1446 138
rect 498 60 544 81
rect 1400 60 1446 81
rect 2272 127 2318 138
rect 2272 60 2318 81
rect 2723 255 2809 453
rect 2902 429 2948 453
rect 2723 209 2742 255
rect 2788 209 2809 255
rect 2723 198 2809 209
rect 2902 255 2948 277
rect 2582 60 2628 81
rect 2902 60 2948 81
rect 0 -60 3024 60
<< via1 >>
rect 1197 554 1249 606
rect 1209 385 1261 393
rect 1209 341 1254 385
rect 1254 341 1261 385
rect 1664 384 1716 393
rect 1664 341 1665 384
rect 1665 341 1711 384
rect 1711 341 1716 384
rect 1786 384 1838 392
rect 1786 340 1831 384
rect 1831 340 1838 384
<< metal2 >>
rect 1183 606 1840 608
rect 1183 554 1197 606
rect 1249 554 1840 606
rect 1183 552 1840 554
rect 1209 395 1265 405
rect 1207 393 1728 395
rect 1207 341 1209 393
rect 1261 341 1664 393
rect 1716 341 1728 393
rect 1207 339 1728 341
rect 1784 392 1840 552
rect 1784 340 1786 392
rect 1838 340 1840 392
rect 1209 329 1265 339
rect 1784 328 1840 340
<< labels >>
flabel metal1 s 0 724 3024 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 3024 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 25 320 172 412 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 797 326 886 586 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel metal1 2723 198 2809 510 0 FreeSans 200 0 0 0 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3024 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 3040 354
string MASKHINTS_PPLUS -16 354 3040 830
<< end >>
