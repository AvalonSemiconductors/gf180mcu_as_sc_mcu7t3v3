magic
tech gf180mcuD
magscale 1 10
timestamp 1764933398
<< nwell >>
rect -86 354 1878 870
<< pwell >>
rect -86 -86 1878 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 940 68 996 268
rect 1104 68 1160 268
rect 1404 68 1460 268
rect 1604 68 1660 268
<< pmos >>
rect 116 440 172 716
rect 372 440 428 716
rect 540 440 596 716
rect 924 440 980 716
rect 1164 440 1220 716
rect 1354 440 1410 716
rect 1604 440 1660 716
<< ndiff >>
rect 28 246 116 268
rect 28 200 41 246
rect 87 200 116 246
rect 28 68 116 200
rect 172 139 276 268
rect 172 93 201 139
rect 247 93 276 139
rect 172 68 276 93
rect 332 246 436 268
rect 332 117 361 246
rect 407 117 436 246
rect 332 68 436 117
rect 492 247 796 268
rect 492 198 737 247
rect 783 198 796 247
rect 492 68 796 198
rect 852 152 940 268
rect 852 106 865 152
rect 911 106 940 152
rect 852 68 940 106
rect 996 127 1104 268
rect 996 81 1029 127
rect 1075 81 1104 127
rect 996 68 1104 81
rect 1160 246 1404 268
rect 1160 198 1299 246
rect 1345 198 1404 246
rect 1160 68 1404 198
rect 1460 239 1604 268
rect 1460 93 1529 239
rect 1575 93 1604 239
rect 1460 68 1604 93
rect 1660 246 1764 268
rect 1660 200 1689 246
rect 1735 200 1764 246
rect 1660 68 1764 200
<< pdiff >>
rect 28 666 116 716
rect 28 488 41 666
rect 87 488 116 666
rect 28 440 116 488
rect 172 686 372 716
rect 172 640 221 686
rect 267 640 372 686
rect 172 440 372 640
rect 428 675 540 716
rect 428 629 457 675
rect 503 629 540 675
rect 428 440 540 629
rect 596 566 684 716
rect 596 468 625 566
rect 671 468 684 566
rect 596 440 684 468
rect 745 663 924 716
rect 745 465 758 663
rect 804 465 924 663
rect 745 440 924 465
rect 980 689 1164 716
rect 980 643 1029 689
rect 1075 643 1164 689
rect 980 440 1164 643
rect 1220 566 1354 716
rect 1220 468 1277 566
rect 1323 468 1354 566
rect 1220 440 1354 468
rect 1410 689 1604 716
rect 1410 643 1519 689
rect 1565 643 1604 689
rect 1410 440 1604 643
rect 1660 666 1764 716
rect 1660 468 1689 666
rect 1735 468 1764 666
rect 1660 440 1764 468
<< ndiffc >>
rect 41 200 87 246
rect 201 93 247 139
rect 361 117 407 246
rect 737 198 783 247
rect 865 106 911 152
rect 1029 81 1075 127
rect 1299 198 1345 246
rect 1529 93 1575 239
rect 1689 200 1735 246
<< pdiffc >>
rect 41 488 87 666
rect 221 640 267 686
rect 457 629 503 675
rect 625 468 671 566
rect 758 465 804 663
rect 1029 643 1075 689
rect 1277 468 1323 566
rect 1519 643 1565 689
rect 1689 468 1735 666
<< polysilicon >>
rect 116 716 172 760
rect 372 716 428 760
rect 540 716 596 760
rect 924 716 980 760
rect 1164 716 1220 760
rect 1354 716 1410 760
rect 1604 716 1660 760
rect 116 396 172 440
rect 372 420 428 440
rect 540 420 596 440
rect 924 420 980 440
rect 1164 420 1220 440
rect 1354 420 1410 440
rect 116 383 193 396
rect 372 384 452 420
rect 116 337 134 383
rect 180 337 193 383
rect 380 377 452 384
rect 116 324 193 337
rect 256 349 328 362
rect 116 268 172 324
rect 256 303 269 349
rect 315 331 328 349
rect 380 331 393 377
rect 439 331 452 377
rect 534 407 606 420
rect 534 361 547 407
rect 593 361 606 407
rect 534 348 606 361
rect 848 407 996 420
rect 848 361 861 407
rect 907 361 996 407
rect 1164 389 1410 420
rect 1604 400 1660 440
rect 1164 384 1221 389
rect 848 348 996 361
rect 315 303 332 331
rect 256 290 332 303
rect 276 268 332 290
rect 380 324 452 331
rect 380 288 492 324
rect 436 268 492 288
rect 940 268 996 348
rect 1044 358 1117 371
rect 1044 312 1057 358
rect 1103 335 1117 358
rect 1208 343 1221 384
rect 1267 384 1410 389
rect 1579 387 1660 400
rect 1267 343 1281 384
rect 1103 312 1160 335
rect 1208 330 1281 343
rect 1456 353 1529 366
rect 1456 335 1469 353
rect 1044 299 1160 312
rect 1104 268 1160 299
rect 1404 307 1469 335
rect 1515 307 1529 353
rect 1579 341 1592 387
rect 1638 341 1660 387
rect 1579 328 1660 341
rect 1404 294 1529 307
rect 1404 268 1460 294
rect 1604 268 1660 328
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 940 24 996 68
rect 1104 24 1160 68
rect 1404 24 1460 68
rect 1604 24 1660 68
<< polycontact >>
rect 134 337 180 383
rect 269 303 315 349
rect 393 331 439 377
rect 547 361 593 407
rect 861 361 907 407
rect 1057 312 1103 358
rect 1221 343 1267 389
rect 1469 307 1515 353
rect 1592 341 1638 387
<< metal1 >>
rect 0 724 1792 844
rect 221 686 267 724
rect 41 666 87 678
rect 1029 689 1075 724
rect 221 629 267 640
rect 446 675 804 678
rect 446 629 457 675
rect 503 663 804 675
rect 503 629 758 663
rect 87 537 576 583
rect 41 267 87 488
rect 134 395 439 490
rect 134 383 180 395
rect 393 377 439 395
rect 134 314 180 337
rect 258 303 269 349
rect 315 303 326 349
rect 530 418 576 537
rect 625 566 671 580
rect 671 468 685 502
rect 625 453 685 468
rect 530 407 593 418
rect 530 361 547 407
rect 530 350 593 361
rect 393 320 439 331
rect 639 318 685 453
rect 258 267 315 303
rect 41 246 315 267
rect 631 272 685 318
rect 1519 689 1565 724
rect 1029 632 1075 643
rect 1137 630 1473 676
rect 1519 632 1565 643
rect 1689 666 1735 678
rect 1137 568 1183 630
rect 1427 583 1473 630
rect 758 313 804 465
rect 872 522 1183 568
rect 1241 566 1381 582
rect 872 407 918 522
rect 850 361 861 407
rect 907 361 918 407
rect 965 430 1195 476
rect 1241 468 1277 566
rect 1323 468 1381 566
rect 1427 537 1689 583
rect 1241 446 1381 468
rect 965 313 1011 430
rect 1149 400 1195 430
rect 1149 389 1267 400
rect 87 220 315 246
rect 361 246 407 258
rect 41 189 87 200
rect 201 139 247 150
rect 631 152 677 272
rect 758 267 1011 313
rect 1057 358 1103 369
rect 1149 343 1221 389
rect 1149 342 1267 343
rect 1221 332 1267 342
rect 758 247 804 267
rect 724 198 737 247
rect 783 198 804 247
rect 1057 221 1103 312
rect 1313 286 1381 446
rect 1427 410 1638 490
rect 1592 387 1638 410
rect 1261 246 1381 286
rect 923 173 1212 221
rect 1261 198 1299 246
rect 1345 198 1381 246
rect 1437 353 1515 364
rect 1437 307 1469 353
rect 1592 330 1638 341
rect 1437 296 1515 307
rect 923 152 971 173
rect 407 117 865 152
rect 361 106 865 117
rect 911 106 971 152
rect 1166 152 1212 173
rect 1437 152 1483 296
rect 201 60 247 93
rect 1018 81 1029 127
rect 1075 81 1086 127
rect 1166 106 1483 152
rect 1529 239 1575 250
rect 1018 60 1086 81
rect 1689 246 1735 468
rect 1689 189 1735 200
rect 1529 60 1575 93
rect 0 -60 1792 60
<< labels >>
flabel metal1 s 0 724 1792 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1792 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 s 134 395 439 490 0 FreeSans 416 0 0 0 EN
port 5 nsew
flabel metal1 s 1427 410 1638 490 0 FreeSans 416 0 0 0 A
port 6 nsew
flabel metal1 s 1313 198 1381 582 0 FreeSans 416 0 0 0 Y
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 1792 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1808 354
string MASKHINTS_PPLUS -16 354 1808 830
<< end >>
