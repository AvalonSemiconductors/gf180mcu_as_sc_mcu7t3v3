magic
tech gf180mcuD
magscale 1 10
timestamp 1751664855
<< nwell >>
rect -86 354 2886 870
<< pwell >>
rect -86 -86 2886 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
rect 1396 68 1452 268
rect 1556 68 1612 268
rect 1716 68 1772 268
rect 1879 68 1935 268
rect 2039 68 2095 268
rect 2199 68 2255 268
rect 2359 68 2415 268
rect 2519 68 2575 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1396 440 1452 716
rect 1556 440 1612 716
rect 1716 440 1772 716
rect 1879 440 1935 716
rect 2039 440 2095 716
rect 2199 440 2255 716
rect 2359 440 2415 716
rect 2519 440 2575 716
<< ndiff >>
rect 28 156 116 268
rect 28 82 41 156
rect 87 82 116 156
rect 28 68 116 82
rect 172 255 276 268
rect 172 209 201 255
rect 247 209 276 255
rect 172 68 276 209
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 255 596 268
rect 492 209 521 255
rect 567 209 596 255
rect 492 68 596 209
rect 652 128 756 268
rect 652 82 681 128
rect 727 82 756 128
rect 652 68 756 82
rect 812 255 916 268
rect 812 209 841 255
rect 887 209 916 255
rect 812 68 916 209
rect 972 127 1076 268
rect 972 81 1001 127
rect 1047 81 1076 127
rect 972 68 1076 81
rect 1132 255 1236 268
rect 1132 209 1161 255
rect 1207 209 1236 255
rect 1132 68 1236 209
rect 1292 127 1396 268
rect 1292 81 1321 127
rect 1367 81 1396 127
rect 1292 68 1396 81
rect 1452 255 1556 268
rect 1452 209 1481 255
rect 1527 209 1556 255
rect 1452 68 1556 209
rect 1612 249 1716 268
rect 1612 81 1641 249
rect 1687 81 1716 249
rect 1612 68 1716 81
rect 1772 255 1879 268
rect 1772 209 1804 255
rect 1850 209 1879 255
rect 1772 68 1879 209
rect 1935 249 2039 268
rect 1935 81 1964 249
rect 2010 81 2039 249
rect 1935 68 2039 81
rect 2095 255 2199 268
rect 2095 209 2124 255
rect 2170 209 2199 255
rect 2095 68 2199 209
rect 2255 249 2359 268
rect 2255 81 2284 249
rect 2330 81 2359 249
rect 2255 68 2359 81
rect 2415 255 2519 268
rect 2415 209 2444 255
rect 2490 209 2519 255
rect 2415 68 2519 209
rect 2575 249 2772 268
rect 2575 81 2604 249
rect 2650 81 2772 249
rect 2575 68 2772 81
<< pdiff >>
rect 28 703 116 716
rect 28 589 41 703
rect 87 589 116 703
rect 28 440 116 589
rect 172 667 276 716
rect 172 472 201 667
rect 247 472 276 667
rect 172 440 276 472
rect 332 701 436 716
rect 332 564 361 701
rect 407 564 436 701
rect 332 440 436 564
rect 492 667 596 716
rect 492 461 521 667
rect 567 461 596 667
rect 492 440 596 461
rect 652 703 756 716
rect 652 565 681 703
rect 727 565 756 703
rect 652 440 756 565
rect 812 667 916 716
rect 812 472 841 667
rect 887 472 916 667
rect 812 440 916 472
rect 972 703 1076 716
rect 972 565 1001 703
rect 1047 565 1076 703
rect 972 440 1076 565
rect 1132 667 1236 716
rect 1132 472 1161 667
rect 1207 472 1236 667
rect 1132 440 1236 472
rect 1292 703 1396 716
rect 1292 564 1321 703
rect 1367 564 1396 703
rect 1292 440 1396 564
rect 1452 667 1556 716
rect 1452 472 1481 667
rect 1527 472 1556 667
rect 1452 440 1556 472
rect 1612 703 1716 716
rect 1612 464 1641 703
rect 1687 464 1716 703
rect 1612 440 1716 464
rect 1772 667 1879 716
rect 1772 453 1804 667
rect 1850 453 1879 667
rect 1772 440 1879 453
rect 1935 703 2039 716
rect 1935 464 1964 703
rect 2010 464 2039 703
rect 1935 440 2039 464
rect 2095 667 2199 716
rect 2095 453 2124 667
rect 2170 453 2199 667
rect 2095 440 2199 453
rect 2255 703 2359 716
rect 2255 464 2284 703
rect 2330 464 2359 703
rect 2255 440 2359 464
rect 2415 667 2519 716
rect 2415 453 2444 667
rect 2490 453 2519 667
rect 2415 440 2519 453
rect 2575 703 2772 716
rect 2575 464 2604 703
rect 2650 464 2772 703
rect 2575 440 2772 464
<< ndiffc >>
rect 41 82 87 156
rect 201 209 247 255
rect 361 81 407 127
rect 521 209 567 255
rect 681 82 727 128
rect 841 209 887 255
rect 1001 81 1047 127
rect 1161 209 1207 255
rect 1321 81 1367 127
rect 1481 209 1527 255
rect 1641 81 1687 249
rect 1804 209 1850 255
rect 1964 81 2010 249
rect 2124 209 2170 255
rect 2284 81 2330 249
rect 2444 209 2490 255
rect 2604 81 2650 249
<< pdiffc >>
rect 41 589 87 703
rect 201 472 247 667
rect 361 564 407 701
rect 521 461 567 667
rect 681 565 727 703
rect 841 472 887 667
rect 1001 565 1047 703
rect 1161 472 1207 667
rect 1321 564 1367 703
rect 1481 472 1527 667
rect 1641 464 1687 703
rect 1804 453 1850 667
rect 1964 464 2010 703
rect 2124 453 2170 667
rect 2284 464 2330 703
rect 2444 453 2490 667
rect 2604 464 2650 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1396 716 1452 760
rect 1556 716 1612 760
rect 1716 716 1772 760
rect 1879 716 1935 760
rect 2039 716 2095 760
rect 2199 716 2255 760
rect 2359 716 2415 760
rect 2519 716 2575 760
rect 116 403 172 440
rect 276 403 332 440
rect 436 403 492 440
rect 596 403 652 440
rect 103 382 652 403
rect 103 336 116 382
rect 629 336 652 382
rect 103 314 652 336
rect 116 268 172 314
rect 276 268 332 314
rect 436 268 492 314
rect 596 268 652 314
rect 756 403 812 440
rect 916 403 972 440
rect 1076 403 1132 440
rect 1236 403 1292 440
rect 1396 403 1452 440
rect 756 381 1452 403
rect 1556 381 1612 440
rect 1716 381 1772 440
rect 1879 381 1935 440
rect 2039 381 2095 440
rect 2199 381 2255 440
rect 2359 381 2415 440
rect 2519 381 2575 440
rect 756 378 2575 381
rect 756 332 769 378
rect 1424 332 2575 378
rect 756 314 1452 332
rect 756 268 812 314
rect 916 268 972 314
rect 1076 268 1132 314
rect 1236 268 1292 314
rect 1396 268 1452 314
rect 1556 268 1612 332
rect 1716 268 1772 332
rect 1879 268 1935 332
rect 2039 268 2095 332
rect 2199 268 2255 332
rect 2359 268 2415 332
rect 2519 268 2575 332
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1396 24 1452 68
rect 1556 24 1612 68
rect 1716 24 1772 68
rect 1879 24 1935 68
rect 2039 24 2095 68
rect 2199 24 2255 68
rect 2359 24 2415 68
rect 2519 24 2575 68
<< polycontact >>
rect 116 336 629 382
rect 769 332 1424 378
<< metal1 >>
rect 0 724 2800 844
rect 41 703 87 724
rect 361 701 407 724
rect 41 570 87 589
rect 201 667 247 678
rect 681 703 727 724
rect 361 553 407 564
rect 521 667 567 678
rect 247 472 521 507
rect 201 461 521 472
rect 1001 703 1047 724
rect 681 554 727 565
rect 841 667 887 678
rect 567 461 721 507
rect 1321 703 1367 724
rect 1001 554 1047 565
rect 1161 667 1207 678
rect 887 472 1161 507
rect 1641 703 1687 724
rect 1321 553 1367 564
rect 1481 667 1527 678
rect 1207 472 1481 507
rect 841 461 1527 472
rect 103 382 629 415
rect 103 336 116 382
rect 103 314 629 336
rect 675 384 721 461
rect 1481 407 1527 461
rect 1964 703 2010 724
rect 1641 453 1687 464
rect 1804 667 1850 678
rect 2284 703 2330 724
rect 1964 453 2010 464
rect 2124 667 2170 678
rect 2604 703 2650 724
rect 2284 453 2330 464
rect 2444 667 2490 678
rect 2604 453 2650 464
rect 1804 407 1850 453
rect 2124 407 2170 453
rect 2444 407 2490 453
rect 675 378 1435 384
rect 675 332 769 378
rect 1424 332 1435 378
rect 675 326 1435 332
rect 675 266 721 326
rect 1481 306 2490 407
rect 1481 266 1527 306
rect 201 255 721 266
rect 247 220 521 255
rect 201 198 247 209
rect 567 220 721 255
rect 841 255 1527 266
rect 521 198 567 209
rect 887 220 1161 255
rect 841 198 887 209
rect 1207 220 1481 255
rect 1161 198 1207 209
rect 1481 198 1527 209
rect 1641 249 1687 260
rect 41 156 87 168
rect 41 60 87 82
rect 361 127 407 142
rect 361 60 407 81
rect 681 128 727 142
rect 681 60 727 82
rect 1001 127 1047 142
rect 1001 60 1047 81
rect 1321 127 1367 142
rect 1321 60 1367 81
rect 1804 255 1850 306
rect 1804 198 1850 209
rect 1964 249 2010 260
rect 1641 60 1687 81
rect 2124 255 2170 306
rect 2124 198 2170 209
rect 2284 249 2330 260
rect 1964 60 2010 81
rect 2444 255 2490 306
rect 2444 198 2490 209
rect 2604 249 2650 260
rect 2284 60 2330 81
rect 2604 60 2650 81
rect 0 -60 2800 60
<< labels >>
flabel metal1 s 0 724 2800 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2800 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 103 314 629 415 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 1481 306 2490 407 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2800 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 2886 354
string MASKHINTS_PPLUS -86 354 2886 870
<< end >>
