magic
tech gf180mcuD
magscale 1 10
timestamp 1753441877
<< nwell >>
rect -86 354 1206 870
<< pwell >>
rect -86 -86 1206 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 724 68 780 268
rect 901 68 957 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 724 440 780 716
rect 901 440 957 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 68 276 268
rect 332 248 436 268
rect 332 202 361 248
rect 407 202 436 248
rect 332 68 436 202
rect 492 127 724 268
rect 492 81 521 127
rect 695 81 724 127
rect 492 68 724 81
rect 780 255 901 268
rect 780 209 826 255
rect 872 209 901 255
rect 780 68 901 209
rect 957 255 1045 268
rect 957 81 986 255
rect 1032 81 1045 255
rect 957 68 1045 81
<< pdiff >>
rect 28 595 116 716
rect 28 549 41 595
rect 87 549 116 595
rect 28 440 116 549
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 595 436 716
rect 332 549 361 595
rect 407 549 436 595
rect 332 440 436 549
rect 492 667 580 716
rect 492 456 521 667
rect 567 456 580 667
rect 492 440 580 456
rect 636 703 724 716
rect 636 453 649 703
rect 695 453 724 703
rect 636 440 724 453
rect 780 665 901 716
rect 780 453 826 665
rect 872 453 901 665
rect 780 440 901 453
rect 957 703 1045 716
rect 957 453 986 703
rect 1032 453 1045 703
rect 957 440 1045 453
<< ndiffc >>
rect 41 81 87 127
rect 361 202 407 248
rect 521 81 695 127
rect 826 209 872 255
rect 986 81 1032 255
<< pdiffc >>
rect 41 549 87 595
rect 201 657 247 703
rect 361 549 407 595
rect 521 456 567 667
rect 649 453 695 703
rect 826 453 872 665
rect 986 453 1032 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 724 716 780 760
rect 901 716 957 760
rect 116 393 172 440
rect 276 393 332 440
rect 436 393 492 440
rect 80 376 172 393
rect 80 330 102 376
rect 148 330 172 376
rect 80 316 172 330
rect 240 377 332 393
rect 240 331 265 377
rect 311 331 332 377
rect 240 316 332 331
rect 400 379 492 393
rect 724 391 780 440
rect 400 333 423 379
rect 469 333 492 379
rect 400 316 492 333
rect 692 377 780 391
rect 901 377 957 440
rect 692 331 714 377
rect 760 331 957 377
rect 692 317 780 331
rect 116 268 172 316
rect 276 268 332 316
rect 436 268 492 316
rect 724 268 780 317
rect 901 268 957 331
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 724 24 780 68
rect 901 24 957 68
<< polycontact >>
rect 102 330 148 376
rect 265 331 311 377
rect 423 333 469 379
rect 714 331 760 377
<< metal1 >>
rect 0 724 1120 844
rect 201 703 247 724
rect 649 703 695 724
rect 201 646 247 657
rect 521 667 567 678
rect 41 595 87 620
rect 361 595 407 609
rect 87 549 361 595
rect 41 533 87 549
rect 361 534 407 549
rect 80 376 172 472
rect 567 456 585 495
rect 521 445 585 456
rect 80 330 102 376
rect 148 330 172 376
rect 80 316 172 330
rect 240 377 332 393
rect 240 331 265 377
rect 311 331 332 377
rect 240 316 332 331
rect 400 379 492 393
rect 400 333 423 379
rect 469 333 492 379
rect 400 316 492 333
rect 539 377 585 445
rect 986 703 1032 724
rect 649 429 695 453
rect 826 665 890 676
rect 872 453 890 665
rect 539 331 714 377
rect 760 331 780 377
rect 539 248 585 331
rect 349 202 361 248
rect 407 202 585 248
rect 826 255 890 453
rect 986 429 1032 453
rect 872 209 890 255
rect 826 198 890 209
rect 986 255 1032 276
rect 41 127 87 138
rect 41 60 87 81
rect 521 127 695 138
rect 521 60 695 81
rect 986 60 1032 81
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 0 724 1120 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1120 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 826 198 890 676 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 80 316 172 472 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 240 316 332 393 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 400 316 492 393 0 FreeSans 200 0 0 0 C
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 1206 354
string MASKHINTS_PPLUS -86 354 1206 870
<< end >>
