magic
tech gf180mcuD
magscale 1 10
timestamp 1751905124
<< nwell >>
rect -86 354 1206 870
<< pwell >>
rect -86 -86 1206 354
<< nmos >>
rect 164 68 220 268
rect 452 68 508 268
rect 612 68 668 268
rect 772 68 828 268
rect 932 68 988 268
<< pmos >>
rect 164 440 220 716
rect 452 440 508 716
rect 612 440 668 716
rect 772 440 828 716
rect 932 440 988 716
<< ndiff >>
rect 72 255 164 268
rect 72 81 89 255
rect 135 81 164 255
rect 72 68 164 81
rect 220 255 308 268
rect 220 209 249 255
rect 295 209 308 255
rect 220 68 308 209
rect 364 218 452 268
rect 364 172 377 218
rect 423 172 452 218
rect 364 68 452 172
rect 508 127 612 268
rect 508 81 537 127
rect 583 81 612 127
rect 508 68 612 81
rect 668 218 772 268
rect 668 172 697 218
rect 743 172 772 218
rect 668 68 772 172
rect 828 255 932 268
rect 828 209 857 255
rect 903 209 932 255
rect 828 68 932 209
rect 988 152 1091 268
rect 988 106 1017 152
rect 1063 106 1091 152
rect 988 68 1091 106
<< pdiff >>
rect 72 703 164 716
rect 72 483 89 703
rect 135 483 164 703
rect 72 440 164 483
rect 220 667 308 716
rect 220 453 249 667
rect 295 453 308 667
rect 220 440 308 453
rect 364 698 452 716
rect 364 483 377 698
rect 423 483 452 698
rect 364 440 452 483
rect 508 621 612 716
rect 508 575 537 621
rect 583 575 612 621
rect 508 440 612 575
rect 668 703 772 716
rect 668 657 697 703
rect 743 657 772 703
rect 668 440 772 657
rect 828 621 932 716
rect 828 575 857 621
rect 903 575 932 621
rect 828 440 932 575
rect 988 703 1092 716
rect 988 657 1018 703
rect 1064 657 1092 703
rect 988 440 1092 657
<< ndiffc >>
rect 89 81 135 255
rect 249 209 295 255
rect 377 172 423 218
rect 537 81 583 127
rect 697 172 743 218
rect 857 209 903 255
rect 1017 106 1063 152
<< pdiffc >>
rect 89 483 135 703
rect 249 453 295 667
rect 377 483 423 698
rect 537 575 583 621
rect 697 657 743 703
rect 857 575 903 621
rect 1018 657 1064 703
<< polysilicon >>
rect 164 716 220 760
rect 452 716 508 760
rect 612 716 668 760
rect 772 716 828 760
rect 932 716 988 760
rect 164 390 220 440
rect 452 404 508 440
rect 134 377 220 390
rect 134 331 147 377
rect 193 331 220 377
rect 134 318 220 331
rect 436 385 508 404
rect 436 339 449 385
rect 495 363 508 385
rect 612 363 668 440
rect 772 403 828 440
rect 932 403 988 440
rect 495 339 668 363
rect 436 323 668 339
rect 164 268 220 318
rect 452 268 508 323
rect 612 268 668 323
rect 762 387 988 403
rect 762 341 775 387
rect 923 341 988 387
rect 762 322 988 341
rect 772 268 828 322
rect 932 268 988 322
rect 164 24 220 68
rect 452 24 508 68
rect 612 24 668 68
rect 772 24 828 68
rect 932 24 988 68
<< polycontact >>
rect 147 331 193 377
rect 449 339 495 385
rect 775 341 923 387
<< metal1 >>
rect 0 724 1120 844
rect 89 703 135 724
rect 377 698 423 724
rect 89 472 135 483
rect 249 667 295 678
rect 697 703 743 724
rect 697 646 743 657
rect 1018 703 1064 724
rect 1018 646 1064 657
rect 537 621 583 632
rect 857 621 903 632
rect 583 575 857 600
rect 903 575 1063 600
rect 537 554 1063 575
rect 377 472 423 483
rect 62 377 202 389
rect 62 331 147 377
rect 193 331 202 377
rect 62 319 202 331
rect 249 383 295 453
rect 436 385 496 404
rect 436 383 449 385
rect 249 339 449 383
rect 495 339 496 385
rect 249 337 496 339
rect 89 255 135 273
rect 249 255 295 337
rect 436 323 496 337
rect 762 387 923 403
rect 762 341 775 387
rect 762 322 923 341
rect 857 264 903 266
rect 969 264 1063 554
rect 857 255 1063 264
rect 249 198 295 209
rect 377 218 743 230
rect 423 184 697 218
rect 377 161 423 172
rect 903 210 1063 255
rect 857 198 903 209
rect 697 152 743 172
rect 89 60 135 81
rect 537 127 583 138
rect 697 106 1017 152
rect 1063 106 1074 152
rect 537 60 583 81
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 0 724 1120 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1120 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 969 210 1063 600 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 762 322 923 403 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 62 319 202 389 0 FreeSans 200 0 0 0 A
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1136 354
string MASKHINTS_PPLUS -16 354 1136 830
<< end >>
