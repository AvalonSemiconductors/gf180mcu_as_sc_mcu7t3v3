magic
tech gf180mcuD
magscale 1 10
timestamp 1753960842
<< nwell >>
rect -86 354 1542 870
<< pwell >>
rect -86 -86 1542 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 189 276 268
rect 172 143 201 189
rect 247 143 276 189
rect 172 68 276 143
rect 332 68 436 268
rect 492 68 596 268
rect 652 127 756 268
rect 652 81 681 127
rect 727 81 756 127
rect 652 68 756 81
rect 812 255 916 268
rect 812 209 841 255
rect 887 209 916 255
rect 812 68 916 209
rect 972 255 1076 268
rect 972 81 1001 255
rect 1047 81 1076 255
rect 972 68 1076 81
rect 1132 255 1236 268
rect 1132 209 1161 255
rect 1207 209 1236 255
rect 1132 68 1236 209
rect 1292 255 1380 268
rect 1292 81 1321 255
rect 1367 81 1380 255
rect 1292 68 1380 81
<< pdiff >>
rect 28 667 116 716
rect 28 453 41 667
rect 87 453 116 667
rect 28 440 116 453
rect 172 600 276 716
rect 172 554 201 600
rect 247 554 276 600
rect 172 440 276 554
rect 332 703 436 716
rect 332 657 361 703
rect 407 657 436 703
rect 332 440 436 657
rect 492 600 596 716
rect 492 554 521 600
rect 567 554 596 600
rect 492 440 596 554
rect 652 703 756 716
rect 652 657 681 703
rect 727 657 756 703
rect 652 440 756 657
rect 812 667 916 716
rect 812 453 841 667
rect 887 453 916 667
rect 812 440 916 453
rect 972 703 1076 716
rect 972 453 1001 703
rect 1047 453 1076 703
rect 972 440 1076 453
rect 1132 667 1236 716
rect 1132 453 1161 667
rect 1207 453 1236 667
rect 1132 440 1236 453
rect 1292 703 1380 716
rect 1292 453 1321 703
rect 1367 453 1380 703
rect 1292 440 1380 453
<< ndiffc >>
rect 41 81 87 127
rect 201 143 247 189
rect 681 81 727 127
rect 841 209 887 255
rect 1001 81 1047 255
rect 1161 209 1207 255
rect 1321 81 1367 255
<< pdiffc >>
rect 41 453 87 667
rect 201 554 247 600
rect 361 657 407 703
rect 521 554 567 600
rect 681 657 727 703
rect 841 453 887 667
rect 1001 453 1047 703
rect 1161 453 1207 667
rect 1321 453 1367 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 116 400 172 440
rect 276 400 332 440
rect 436 400 492 440
rect 596 400 652 440
rect 756 400 812 440
rect 116 380 198 400
rect 116 334 139 380
rect 185 334 198 380
rect 116 317 198 334
rect 276 382 358 400
rect 276 336 290 382
rect 336 336 358 382
rect 276 317 358 336
rect 436 378 518 400
rect 436 332 453 378
rect 499 332 518 378
rect 436 317 518 332
rect 596 383 678 400
rect 596 337 613 383
rect 659 337 678 383
rect 596 317 678 337
rect 736 383 812 400
rect 916 383 972 440
rect 1076 383 1132 440
rect 1236 383 1292 440
rect 736 337 749 383
rect 795 337 1292 383
rect 736 317 812 337
rect 116 268 172 317
rect 276 268 332 317
rect 436 268 492 317
rect 596 268 652 317
rect 756 268 812 317
rect 916 268 972 337
rect 1076 268 1132 337
rect 1236 268 1292 337
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
<< polycontact >>
rect 139 334 185 380
rect 290 336 336 382
rect 453 332 499 378
rect 613 337 659 383
rect 749 337 795 383
<< metal1 >>
rect 0 724 1456 844
rect 361 703 407 724
rect 41 667 87 678
rect 361 646 407 657
rect 681 703 727 724
rect 1001 703 1047 724
rect 681 646 727 657
rect 841 667 909 678
rect 190 554 201 600
rect 247 554 521 600
rect 567 554 580 600
rect 41 230 87 453
rect 133 380 217 487
rect 133 334 139 380
rect 185 334 217 380
rect 133 317 217 334
rect 276 382 360 487
rect 887 453 909 667
rect 276 336 290 382
rect 336 336 360 382
rect 276 317 360 336
rect 436 378 520 400
rect 436 332 453 378
rect 499 332 520 378
rect 436 230 520 332
rect 596 383 664 421
rect 749 383 795 394
rect 596 337 613 383
rect 659 337 664 383
rect 596 317 664 337
rect 726 337 749 383
rect 726 326 795 337
rect 841 382 909 453
rect 1321 703 1367 724
rect 1001 436 1047 453
rect 1161 667 1229 678
rect 1207 453 1229 667
rect 1161 382 1229 453
rect 1321 436 1367 453
rect 841 336 1229 382
rect 726 230 772 326
rect 41 189 247 230
rect 41 184 201 189
rect 589 184 772 230
rect 841 255 909 336
rect 887 209 909 255
rect 841 198 909 209
rect 1001 255 1047 274
rect 589 152 635 184
rect 247 143 635 152
rect 41 127 87 138
rect 201 106 635 143
rect 681 127 727 138
rect 41 60 87 81
rect 681 60 727 81
rect 1161 255 1229 336
rect 1207 209 1229 255
rect 1161 198 1229 209
rect 1321 255 1367 274
rect 1001 60 1047 81
rect 1321 60 1367 81
rect 0 -60 1456 60
<< labels >>
flabel metal1 s 0 724 1456 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1456 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 133 317 217 487 0 FreeSans 200 0 0 0 D
port 5 nsew signal input
flabel metal1 276 317 360 487 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 436 230 520 400 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 596 317 664 421 0 FreeSans 200 0 0 0 C
port 8 nsew signal input
flabel metal1 841 198 909 678 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel metal1 1161 198 1229 678 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 1472 354
string MASKHINTS_PPLUS -16 354 1472 830
<< end >>
