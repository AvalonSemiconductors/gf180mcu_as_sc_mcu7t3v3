magic
tech gf180mcuD
magscale 1 10
timestamp 1758890550
<< nwell >>
rect -86 354 310 870
<< pwell >>
rect -86 -86 310 354
<< psubdiff >>
rect 56 245 168 258
rect 56 70 86 245
rect 132 70 168 245
rect 56 56 168 70
<< nsubdiff >>
rect 72 665 152 712
rect 72 431 86 665
rect 132 431 152 665
rect 72 384 152 431
<< psubdiffcont >>
rect 86 70 132 245
<< nsubdiffcont >>
rect 86 431 132 665
<< metal1 >>
rect 0 724 224 844
rect 75 665 143 724
rect 75 431 86 665
rect 132 431 143 665
rect 75 386 143 431
rect 75 245 143 302
rect 75 70 86 245
rect 132 70 143 245
rect 75 60 143 70
rect 0 -60 224 60
<< labels >>
flabel metal1 s 0 724 224 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 224 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 784
string LEFclass CORE WELLTAP
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 310 354
string MASKHINTS_PPLUS -86 354 310 870
<< end >>
