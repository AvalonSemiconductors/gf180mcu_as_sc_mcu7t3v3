magic
tech gf180mcuD
magscale 1 10
timestamp 1753182340
<< nwell >>
rect -86 354 1318 870
<< pwell >>
rect -86 -86 1318 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 884 68 940 268
rect 1044 68 1100 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 884 440 940 716
rect 1044 440 1100 716
<< ndiff >>
rect 28 255 116 268
rect 28 81 41 255
rect 87 81 116 255
rect 28 68 116 81
rect 172 224 276 268
rect 172 178 201 224
rect 247 178 276 224
rect 172 68 276 178
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 223 596 268
rect 492 177 521 223
rect 567 177 596 223
rect 492 68 596 177
rect 652 132 884 268
rect 652 86 681 132
rect 855 86 884 132
rect 652 68 884 86
rect 940 251 1044 268
rect 940 205 969 251
rect 1015 205 1044 251
rect 940 68 1044 205
rect 1100 255 1190 268
rect 1100 81 1129 255
rect 1175 81 1190 255
rect 1100 68 1190 81
<< pdiff >>
rect 28 575 116 716
rect 28 529 41 575
rect 87 529 116 575
rect 28 440 116 529
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 628 436 716
rect 332 582 361 628
rect 407 582 436 628
rect 332 440 436 582
rect 492 575 596 716
rect 492 529 521 575
rect 567 529 596 575
rect 492 440 596 529
rect 652 671 740 716
rect 652 625 681 671
rect 727 625 740 671
rect 652 440 740 625
rect 796 625 884 716
rect 796 579 809 625
rect 855 579 884 625
rect 796 440 884 579
rect 940 550 1044 716
rect 940 453 969 550
rect 1015 453 1044 550
rect 940 440 1044 453
rect 1100 655 1190 716
rect 1100 453 1129 655
rect 1175 453 1190 655
rect 1100 440 1190 453
<< ndiffc >>
rect 41 81 87 255
rect 201 178 247 224
rect 361 81 407 127
rect 521 177 567 223
rect 681 86 855 132
rect 969 205 1015 251
rect 1129 81 1175 255
<< pdiffc >>
rect 41 529 87 575
rect 201 657 247 703
rect 361 582 407 628
rect 521 529 567 575
rect 681 625 727 671
rect 809 579 855 625
rect 969 453 1015 550
rect 1129 453 1175 655
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 884 716 940 760
rect 1044 716 1100 760
rect 116 394 172 440
rect 276 394 332 440
rect 75 380 332 394
rect 436 391 492 440
rect 596 391 652 440
rect 884 394 940 440
rect 75 334 88 380
rect 285 334 332 380
rect 75 317 332 334
rect 116 268 172 317
rect 276 268 332 317
rect 395 375 652 391
rect 395 329 408 375
rect 639 329 652 375
rect 395 314 652 329
rect 836 378 940 394
rect 1044 378 1100 440
rect 836 332 850 378
rect 896 332 1100 378
rect 836 317 940 332
rect 436 268 492 314
rect 596 268 652 314
rect 884 268 940 317
rect 1044 268 1100 332
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 884 24 940 68
rect 1044 24 1100 68
<< polycontact >>
rect 88 334 285 380
rect 408 329 639 375
rect 850 332 896 378
<< metal1 >>
rect 0 724 1232 844
rect 201 703 247 724
rect 201 646 247 657
rect 361 628 681 671
rect 41 575 87 586
rect 407 625 681 628
rect 727 625 738 671
rect 809 655 1175 666
rect 809 625 1129 655
rect 361 575 407 582
rect 855 620 1129 625
rect 809 575 855 579
rect 87 530 407 575
rect 87 529 382 530
rect 510 529 521 575
rect 567 529 855 575
rect 969 550 1036 561
rect 41 518 87 529
rect 75 380 285 394
rect 75 334 88 380
rect 75 317 285 334
rect 395 375 652 391
rect 395 329 408 375
rect 639 329 652 375
rect 395 314 652 329
rect 836 378 916 483
rect 836 332 850 378
rect 896 332 916 378
rect 836 317 916 332
rect 1015 453 1036 550
rect 41 255 87 271
rect 969 251 1036 453
rect 1129 425 1175 453
rect 201 224 969 251
rect 247 223 969 224
rect 247 205 521 223
rect 201 167 247 178
rect 567 205 969 223
rect 1015 205 1036 251
rect 1129 255 1175 274
rect 521 166 567 177
rect 41 60 87 81
rect 361 127 407 143
rect 361 60 407 81
rect 681 132 855 143
rect 681 60 855 86
rect 1129 60 1175 81
rect 0 -60 1232 60
<< labels >>
flabel metal1 s 0 724 1232 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1232 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 75 317 285 394 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 395 314 652 391 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 836 317 916 483 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 969 205 1036 550 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1232 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
string MASKHINTS_NPLUS -86 -86 1318 354
string MASKHINTS_PPLUS -86 354 1318 870
<< end >>
