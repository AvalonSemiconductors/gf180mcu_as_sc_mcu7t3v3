.option method=key

.param
+  sw_stat_global = 0
+  sw_stat_mismatch = 0
+ mc_skew = 3
+ res_mc_skew = 3
+ cap_mc_skew = 3
+  fnoicor = 0

.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.option wnflag=1

.include ./gf180mcu_extra__dffm2_2.spice

VDD VDD 0 3.3V
VSS VSS 0 0V

R1111 VNW GND 0
R1121 VPW VDD 0
R1131 GND VSS 0

Va D0 GND PULSE( 0 3.3 20ns 0.1ns 0.1ns 10ns 50ns )
Vb CLK GND PULSE( 0 3.3 5ns 0.1ns 0.1ns 10ns 20ns )

.tran 1n 60n

.control
run
plot v(CLK)+4 v(D0)+2 v(Q0)
.endc
.end
